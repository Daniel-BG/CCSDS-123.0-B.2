----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02.03.2021 10:35:20
-- Design Name: 
-- Module Name: constants - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.ccsds_math_functions.all;

package ccsds_constants is
	constant TEST_GEN_ENABLE: boolean := false;

	--IMAGE CONSTANTS
	type relocation_mode_t is (VERTICAL_TO_DIAGONAL, DIAGONAL_TO_VERTICAL); 
	
	--OTHER CONSTANTS
	constant STDLV_ONE: std_logic_vector(0 downto 0) := "1";
	constant STDLV_ZERO: std_logic_vector(0 downto 0) := "0";
	
	--FIXED CONSTANTS
	constant CONST_TINC_MIN				: integer := 4;
	constant CONST_TINC_MAX				: integer := 11;
	constant CONST_TINC_BITS 			: integer := 4;
	constant CONST_VMIN					: integer := -6;
	constant CONST_VMAX					: integer := 9;
	constant CONST_VMINMAX_BITS 		: integer := 5;
	constant CONST_WEO_MIN				: integer := -6;
	constant CONST_WEO_MAX				: integer := 5;
	constant CONST_WEO_BITS 			: integer := 4;
	constant CONST_MAX_RES_VAL 			: integer := 4;
	constant CONST_DATA_WIDTH_MAX		: integer := 32;
	constant CONST_DATA_WIDTH_MIN		: integer := 2;
	constant CONST_OMEGA_WIDTH_MAX		: integer := 19;
	constant CONST_OMEGA_WIDTH_MIN		: integer := 4;
	constant CONST_WUSE_BITS 			: integer := 7;

	--CONSTANTS THAT CAN ALTER RESOURCE USE
	constant CONST_MAX_DATA_WIDTH		: integer := 16;				--maximum allowed bits for inputs (Can be set lower through cfg ports)
	constant CONST_MAX_OMEGA			: integer := 19;				--maximum allowed bits for weights (Can be set lower through cfg ports)
	constant CONST_MIN_OMEGA			: integer := 4;
	constant CONST_MAX_P				: integer := 3;					--maximum allowed bits for previous bands used in prediction
	constant CONST_MAX_BANDS			: integer := 32;				--maximum allowed size in the z direction (Can be set lower through cfg ports)
	constant CONST_MAX_LINES			: integer := 64;				--maximum allowed size in the y direction (Can be set lower through cfg ports)
	constant CONST_MAX_SAMPLES			: integer := 128; 				--maximum allowed size in the x direction (Can be set lower through cfg ports)
	
	--DERIVED CONSTANTS
	constant CONST_MAX_SAMPLES_PER_BAND	: integer := CONST_MAX_SAMPLES * CONST_MAX_LINES;
	
	constant CONST_MAX_X_VALUE			: integer := CONST_MAX_SAMPLES - 1;	--maximum allowed size in the x direction (Can be set lower through cfg ports)
	constant CONST_MAX_Y_VALUE			: integer := CONST_MAX_LINES - 1;	--maximum allowed size in the y direction (Can be set lower through cfg ports)
	constant CONST_MAX_Z_VALUE			: integer := CONST_MAX_BANDS - 1;  	--maximum allowed size in the z direction (Can be set lower through cfg ports)
	constant CONST_MAX_T_VALUE			: integer := CONST_MAX_SAMPLES_PER_BAND - 1;
	
	constant CONST_ABS_ERR_BITS 		: integer := MIN(CONST_MAX_DATA_WIDTH - 1, 16); 
	constant CONST_REL_ERR_BITS 		: integer := MIN(CONST_MAX_DATA_WIDTH - 1, 16); 
	
	constant CONST_MAX_WEIGHT_BITS		: integer := CONST_MAX_OMEGA + 3;
	constant CONST_MAX_C				: integer := CONST_MAX_P + 3; --number of previous bands plus 3 (full pred mode)
	constant CONST_MAX_OMEGA_WIDTH_BITS	: integer := BITS(CONST_MAX_OMEGA);		
	constant CONST_MAX_DATA_WIDTH_BITS	: integer := BITS(CONST_MAX_DATA_WIDTH);	
	constant CONST_MAX_P_WIDTH_BITS  	: integer := BITS(CONST_MAX_P);
	constant CONST_MAX_C_BITS			: integer := BITS(CONST_MAX_C);
	
	constant CONST_MAX_X_VALUE_BITS		: integer := BITS(CONST_MAX_X_VALUE);
	constant CONST_MAX_Y_VALUE_BITS		: integer := BITS(CONST_MAX_Y_VALUE);
	constant CONST_MAX_Z_VALUE_BITS		: integer := BITS(CONST_MAX_Z_VALUE);
	constant CONST_MAX_T_VALUE_BITS		: integer := BITS(CONST_MAX_T_VALUE);
	
	constant CONST_MAX_BANDS_BITS		: integer := BITS(CONST_MAX_BANDS);
	constant CONST_MAX_LINES_BITS		: integer := BITS(CONST_MAX_LINES);
	constant CONST_MAX_SAMPLES_BITS		: integer := BITS(CONST_MAX_SAMPLES);
	
	constant CONST_CQBC_BITS			: integer := CONST_MAX_DATA_WIDTH;
	constant CONST_QI_BITS				: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_LSUM_BITS			: integer := CONST_MAX_DATA_WIDTH + 2;
	constant CONST_LDIF_BITS			: integer := CONST_MAX_DATA_WIDTH + 3;
	constant CONST_DRSR_BITS 			: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_DRPSV_BITS 			: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_DRPE_BITS 			: integer := CONST_MAX_DATA_WIDTH + 2;
	constant CONST_PR_BITS 				: integer := CONST_MAX_DATA_WIDTH + 1;
	
	constant CONST_MEV_BITS 			: integer := MAX(CONST_ABS_ERR_BITS, CONST_REL_ERR_BITS);
	constant CONST_PCLD_BITS 			: integer := CONST_MAX_WEIGHT_BITS + CONST_MAX_DATA_WIDTH + BITS(8*CONST_MAX_P + 19);
	constant CONST_HRPSV_BITS			: integer := CONST_MAX_OMEGA + 2 + CONST_MAX_DATA_WIDTH;
	
	constant CONST_RES_BITS				: integer := BITS(CONST_MAX_RES_VAL);
	constant CONST_DAMPING_BITS			: integer := CONST_MAX_RES_VAL;
	constant CONST_OFFSET_BITS			: integer := CONST_MAX_RES_VAL;
	
	constant CONST_DIFFVEC_BITS 		: integer := CONST_MAX_C * CONST_LDIF_BITS;
	constant CONST_CLDVEC_BITS 			: integer := CONST_MAX_P * CONST_LDIF_BITS;
	constant CONST_DIRDIFFVEC_BITS		: integer := 3 * CONST_LDIF_BITS;
	constant CONST_WEIGHTVEC_BITS		: integer := CONST_MAX_C * CONST_MAX_WEIGHT_BITS;
	
	constant CONST_W_UPDATE_BITS		: integer := CONST_LDIF_BITS - CONST_VMIN - CONST_WEO_MIN - CONST_DATA_WIDTH_MIN + CONST_OMEGA_WIDTH_MAX; --should be 64
	
	constant CONST_THETA_BITS			: integer := CONST_MAX_DATA_WIDTH;
	constant CONST_MQI_BITS				: integer := CONST_MAX_DATA_WIDTH;
	
	--ENCODER OUTPUT CONSTANTS
	constant CONST_OUTPUT_CODE_LENGTH 	: integer := 64;
	constant CONST_OUTPUT_CODE_LENGTH_BITS: integer := 7;
	
	--ENCODER CONSTANTS
	constant CONST_MIN_GAMMA_ZERO		: integer := 1;
	constant CONST_MAX_GAMMA_ZERO		: integer := 8;
	constant CONST_MAX_GAMMA_STAR		: integer := 11;
	constant CONST_MAX_GAMMA_STAR_BITS	: integer := BITS(CONST_MAX_GAMMA_STAR);
	constant CONST_MAX_COUNTER_BITS 	: integer := CONST_MAX_GAMMA_STAR;
	constant CONST_MAX_ACC_BITS			: integer := CONST_MAX_GAMMA_STAR + CONST_MAX_DATA_WIDTH;
	constant CONST_MAX_HR_ACC_BITS		: integer := CONST_MAX_ACC_BITS + 2;
	constant CONST_MAX_K				: integer := CONST_MAX_DATA_WIDTH - 2;
	constant CONST_MAX_K_BITS			: integer := BITS(CONST_MAX_K);
	constant CONST_U_MAX_MIN			: integer := 8;
	constant CONST_U_MAX_MAX			: integer := 32;
	constant CONST_U_MAX_BITS			: integer := BITS(CONST_U_MAX_MAX);
	
	constant CONST_MAX_CODE_LENGTH		: integer := CONST_U_MAX_MAX + CONST_MAX_DATA_WIDTH;
	constant CONST_MAX_CODE_LENGTH_BITS : integer := BITS(CONST_MAX_CODE_LENGTH);
	
	--HYBRID ENCODER SPECIFIC CONSTANTS
	constant CONST_LE_TABLE_COUNT: integer := 16;
	constant CONST_CODE_INDEX_BITS: integer := bits(CONST_LE_TABLE_COUNT - 1);
	
	constant CONST_MAX_THRESHOLD_VALUE_BITS : integer := 19;
	subtype threshold_value_t is std_logic_vector (CONST_MAX_THRESHOLD_VALUE_BITS - 1 downto 0);
    type threshold_table_t is array (0 to CONST_LE_TABLE_COUNT - 1) of threshold_value_t;

    constant CONST_THRESHOLD_TABLE : threshold_table_t := (
		"100" & x"A0E8",
		"011" & x"707C",
		"010" & x"8C43",
		"001" & x"F6A0",
		"001" & x"756D",
		"001" & x"1026",
		"000" & x"C5F6",
		"000" & x"8852",
		"000" & x"5B23",
		"000" & x"3A57",
		"000" & x"2442",
		"000" & x"1586",
		"000" & x"0C7B",
		"000" & x"0788",
		"000" & x"0458",
		"000" & x"0198"
	);
	
	constant CONST_INPUT_SYMBOL_AMOUNT: integer := 15;
	constant CONST_INPUT_SYMBOL_BITS: integer := bits(CONST_INPUT_SYMBOL_AMOUNT - 1);
	constant CONST_INPUT_SYMBOL_X	 : std_logic_vector := std_logic_vector(to_unsigned(13, CONST_INPUT_SYMBOL_BITS)); --"1101";
	constant CONST_INPUT_SYMBOL_FLUSH: std_logic_vector := std_logic_vector(to_unsigned(14, CONST_INPUT_SYMBOL_BITS)); --"1110";
	
	type input_symbol_limit_t is array (0 to CONST_LE_TABLE_COUNT - 1) of std_logic_vector(CONST_INPUT_SYMBOL_BITS - 1 downto 0);
	constant CONST_INPUT_SYMBOL_LIMIT : input_symbol_limit_t := (
		x"C", x"A", x"8", x"6",
		x"6", x"4", x"4", x"4",
		x"2", x"2", x"2", x"2",
		x"2", x"2", x"2", x"0"		
	);
	
	constant CONST_CODEWORD_BITS: integer := 21;
	constant CONST_CODEWORD_LENGTH_BITS: integer := 5;
	
	constant CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT: integer := 688;
	constant CONST_LOW_ENTROPY_CODING_TABLE_ADDRESS_BITS: integer := bits(CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT);
	
	constant CONST_LOW_ENTROPY_TABLE_ENTRY_BITS: integer := 40;

	type table_rom_t_v2 is array(0 to CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT*16 - 1) of std_logic_vector(CONST_LOW_ENTROPY_TABLE_ENTRY_BITS - 1 downto 0);
	constant CONST_LOW_ENTROPY_CODING_TABLE_V2: table_rom_t_v2 := (
		x"c000000010",x"4180000000",x"4180001000",x"4180000800",x"c000000011",x"4200001800",x"4200003800",x"c000000012",x"c000000013",x"4280000400",x"4280004400",x"4300001400",x"4300009400",x"4280002400",x"7080000000",x"3000000000",
		x"c000000014",x"c000000015",x"c000000016",x"4180000001",x"4180001001",x"4200000801",x"4200002801",x"4280001801",x"4280005801",x"4300003401",x"c000000017",x"3000000000",x"3000000000",x"430000b401",x"7080000000",x"3000000000",
		x"4100000002",x"c000000018",x"c000000019",x"4180000802",x"4180001802",x"c00000001a",x"c00000001b",x"4300006402",x"430000e402",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4300001402",x"7080000000",x"3000000000",
		x"c00000001c",x"4100000003",x"c00000001d",x"c00000001e",x"c00000001f",x"4280003803",x"c000000020",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4300001403",x"7080000000",x"3000000000",
		x"c000000021",x"4100000004",x"4100000804",x"4200000404",x"4200002404",x"4380004c04",x"4380014c04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4400009c04",x"7080000000",x"3000000000",
		x"4080000005",x"4100000405",x"c000000022",x"4280000c05",x"4280004c05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4380006c05",x"7080000000",x"3000000000",
		x"c000000023",x"c000000024",x"c000000025",x"c000000026",x"4380002c06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001bc06",x"7100000000",x"3000000000",
		x"c000000027",x"c000000028",x"4180000407",x"c000000029",x"448003bc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"450006fc07",x"7080000000",x"3000000000",
		x"c00000002a",x"c00000002b",x"c00000002c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001bc08",x"7100000000",x"3000000000",
		x"c00000002d",x"4200000809",x"4200002809",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4500017c09",x"7180000000",x"3000000000",
		x"c00000002e",x"c00000002f",x"428000040a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460017fc0a",x"7180000000",x"3000000000",
		x"c000000030",x"428000040b",x"c000000031",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47002ffc0b",x"7200000000",x"3000000000",
		x"c000000032",x"430000040c",x"430000840c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47806ffc0c",x"7200000000",x"3000000000",
		x"c000000033",x"c000000034",x"438000040d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47800ffc0d",x"7280000000",x"3000000000",
		x"c000000035",x"440000040e",x"440002040e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48000ffc0e",x"7300000000",x"3000000000",
		x"c000000036",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000040f",x"7400000000",x"3000000000",
		x"4280006400",x"c000000037",x"c000000038",x"4300005400",x"430000d400",x"4300003400",x"430000b400",x"4380004c00",x"4380014c00",x"440000ec00",x"440002ec00",x"4480003c00",x"4480043c00",x"440001ec00",x"7100000400",x"3000000000",
		x"4300007400",x"430000f400",x"4300000c00",x"4300008c00",x"c000000039",x"438000cc00",x"438001cc00",x"440003ec00",x"4400001c00",x"4480023c00",x"4480063c00",x"4480013c00",x"4480053c00",x"4400021c00",x"7180000c00",x"3000000000",
		x"4380002c00",x"4380012c00",x"438000ac00",x"4400011c00",x"4400031c00",x"4400009c00",x"4400029c00",x"4480033c00",x"4480073c00",x"4500057c00",x"45000d7c00",x"458001fc00",x"458011fc00",x"4500037c00",x"7280001c00",x"3000000000",
		x"438001ac00",x"4380006c00",x"4380016c00",x"4400019c00",x"4400039c00",x"4400005c00",x"4400025c00",x"448000bc00",x"448004bc00",x"45000b7c00",x"4500077c00",x"458009fc00",x"458019fc00",x"45000f7c00",x"7280005c00",x"3000000000",
		x"c00000003a",x"4280003801",x"4280007801",x"c00000003b",x"c00000003c",x"4300007401",x"430000f401",x"4380004c01",x"4380014c01",x"4480039c01",x"4480079c01",x"3000000000",x"3000000000",x"440000ac01",x"7180000400",x"3000000000",
		x"4280000401",x"4280004401",x"4280002401",x"c00000003d",x"4300000c01",x"c00000003e",x"c00000003f",x"440002ac01",x"440001ac01",x"4480005c01",x"4480045c01",x"3000000000",x"3000000000",x"4480025c01",x"7180001400",x"3000000000",
		x"4280006401",x"4280001401",x"4280005401",x"c000000040",x"4300008c01",x"c000000041",x"438000cc01",x"440003ac01",x"4400006c01",x"4480065c01",x"4480015c01",x"3000000000",x"3000000000",x"4480055c01",x"7180000c00",x"3000000000",
		x"4480035c01",x"4480075c01",x"448000dc01",x"450007bc01",x"45000fbc01",x"4500007c01",x"4500087c01",x"458008fc01",x"460005fc01",x"468037fc01",x"468077fc01",x"3000000000",x"3000000000",x"460025fc01",x"7380007c00",x"3000000000",
		x"4200000402",x"c000000042",x"c000000043",x"c000000044",x"c000000045",x"438000d402",x"438001d402",x"440001ac02",x"448003dc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007dc02",x"7180000400",x"3000000000",
		x"c000000046",x"c000000047",x"4280002402",x"c000000048",x"c000000049",x"4380003402",x"4380013402",x"440003ac02",x"4480003c02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480043c02",x"7180001400",x"3000000000",
		x"4300009402",x"438000b402",x"438001b402",x"4400006c02",x"4400026c02",x"4480023c02",x"4480063c02",x"458002fc02",x"458012fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45800afc02",x"7280000c00",x"3000000000",
		x"4380007402",x"4380017402",x"438000f402",x"4400016c02",x"4400036c02",x"4480013c02",x"4480053c02",x"45801afc02",x"458006fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458016fc02",x"7280004c00",x"3000000000",
		x"c00000004a",x"4200000803",x"4200002803",x"4280007803",x"4280000403",x"438000b403",x"438001b403",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"440001ac03",x"7180000400",x"3000000000",
		x"4200001803",x"c00000004b",x"c00000004c",x"c00000004d",x"4300009403",x"440003ac03",x"4400006c03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4400026c03",x"7180001400",x"3000000000",
		x"4280004403",x"c00000004e",x"c00000004f",x"4380007403",x"4380017403",x"448001dc03",x"448005dc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003dc03",x"7200000c00",x"3000000000",
		x"4280002403",x"c000000050",x"4300005403",x"438000f403",x"438001f403",x"448007dc03",x"4480003c03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4500037c03",x"7280001c00",x"3000000000",
		x"4380000c03",x"4400016c03",x"4400036c03",x"4480043c03",x"4480023c03",x"45800afc03",x"45801afc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46000bfc03",x"7380003c00",x"3000000000",
		x"c000000051",x"c000000052",x"c000000053",x"c000000054",x"c000000055",x"4400029c04",x"4400019c04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003bc04",x"7100000400",x"3000000000",
		x"c000000056",x"c000000057",x"c000000058",x"4380016c05",x"c000000059",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002dc05",x"7180000400",x"3000000000",
		x"c00000005a",x"4180000006",x"c00000005b",x"4380012c06",x"438000ac06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005bc06",x"7100000800",x"3000000000",
		x"4180001006",x"c00000005c",x"4280002406",x"448003bc06",x"448007bc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458006fc06",x"7200001400",x"3000000000",
		x"c00000005d",x"4280006406",x"4280001406",x"4480007c06",x"4480047c06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458016fc06",x"7200003400",x"3000000000",
		x"438001ac06",x"4480027c06",x"4480067c06",x"468017fc06",x"468057fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780fffc06",x"740001fc00",x"3000000000",
		x"4080000007",x"c00000005e",x"c00000005f",x"448007bc07",x"4480007c07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458009fc07",x"7100000400",x"3000000000",
		x"c000000060",x"c000000061",x"4300002c07",x"458019fc07",x"458005fc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46800ffc07",x"7200000c00",x"3000000000",
		x"4480047c07",x"458015fc07",x"45800dfc07",x"48007ffc07",x"4882fffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4907fffc07",x"748003fc00",x"3000000000",
		x"c000000062",x"c000000063",x"4200001008",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005bc08",x"7180000800",x"3000000000",
		x"c000000064",x"c000000065",x"4380006c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460007fc08",x"7300001c00",x"3000000000",
		x"c000000066",x"c000000067",x"4380016c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460027fc08",x"7300009c00",x"3000000000",
		x"c000000068",x"4200001809",x"c000000069",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458003fc09",x"7180001000",x"3000000000",
		x"c00000006a",x"c00000006b",x"428000440a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460037fc0a",x"7180001000",x"3000000000",
		x"c00000006c",x"448000bc0a",x"450006bc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48807ffc0a",x"7400003c00",x"3000000000",
		x"c00000006d",x"c00000006e",x"c00000006f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700affc0b",x"7200002000",x"3000000000",
		x"c000000070",x"4580017c0b",x"4580117c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a0dfffc0b",x"7500037c00",x"3000000000",
		x"c000000071",x"430000440c",x"c000000072",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47816ffc0c",x"7200002000",x"3000000000",
		x"c000000073",x"438001040d",x"438000840d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47810ffc0d",x"7280004000",x"3000000000",
		x"c000000074",x"460007fc0d",x"460027fc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4907fffc0d",x"740001fc00",x"3000000000",
		x"c000000075",x"440001040e",x"440003040e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48020ffc0e",x"7300008000",x"3000000000",
		x"c000000076",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004040f",x"7400020000",x"3000000000",
		x"4400015c00",x"4400035c00",x"440000dc00",x"448002bc00",x"448006bc00",x"448001bc00",x"448005bc00",x"450000fc00",x"450008fc00",x"458005fc00",x"458015fc00",x"460007fc00",x"460027fc00",x"45800dfc00",x"7280003c00",x"3000000000",
		x"440002dc00",x"440001dc00",x"440003dc00",x"448003bc00",x"448007bc00",x"4480007c00",x"4480047c00",x"450004fc00",x"45000cfc00",x"45801dfc00",x"458003fc00",x"460017fc00",x"460037fc00",x"458013fc00",x"7300007c00",x"3000000000",
		x"4480027c00",x"4480067c00",x"4480017c00",x"450002fc00",x"45000afc00",x"450006fc00",x"45000efc00",x"45800bfc00",x"45801bfc00",x"46000ffc00",x"46002ffc00",x"46803ffc00",x"46807ffc00",x"46001ffc00",x"730000fc00",x"3000000000",
		x"438001cc01",x"4380002c01",x"4380012c01",x"4400026c01",x"4400016c01",x"448004dc01",x"448002dc01",x"4500047c01",x"45000c7c01",x"458018fc01",x"458004fc01",x"3000000000",x"3000000000",x"458014fc01",x"7280001c00",x"3000000000",
		x"4400036c01",x"440000ec01",x"440002ec01",x"448006dc01",x"448001dc01",x"448005dc01",x"448003dc01",x"4500027c01",x"45800cfc01",x"460015fc01",x"460035fc01",x"3000000000",x"3000000000",x"45801cfc01",x"7300005c00",x"3000000000",
		x"440001ec01",x"440003ec01",x"4400001c01",x"448007dc01",x"4480003c01",x"4480043c01",x"45000a7c01",x"458002fc01",x"458012fc01",x"46000dfc01",x"46002dfc01",x"3000000000",x"3000000000",x"45800afc01",x"730000dc00",x"3000000000",
		x"4400021c01",x"4400011c01",x"4400031c01",x"4480023c01",x"4480063c01",x"4500067c01",x"45000e7c01",x"45801afc01",x"458006fc01",x"46001dfc01",x"46003dfc01",x"3000000000",x"3000000000",x"460003fc01",x"7300003c00",x"3000000000",
		x"4480013c01",x"4480053c01",x"4480033c01",x"4500017c01",x"4500097c01",x"4500057c01",x"458016fc01",x"460023fc01",x"460013fc01",x"46800ffc01",x"46804ffc01",x"3000000000",x"3000000000",x"460033fc01",x"7380017c00",x"3000000000",
		x"4480073c01",x"448000bc01",x"448004bc01",x"45000d7c01",x"4500037c01",x"45800efc01",x"45801efc01",x"46000bfc01",x"46002bfc01",x"46802ffc01",x"46806ffc01",x"3000000000",x"3000000000",x"46801ffc01",x"738000fc00",x"3000000000",
		x"4400009c01",x"4400029c01",x"4400019c01",x"448002bc01",x"448006bc01",x"45000b7c01",x"4500077c01",x"458001fc01",x"458011fc01",x"46001bfc01",x"46003bfc01",x"3000000000",x"3000000000",x"460007fc01",x"730000bc00",x"3000000000",
		x"448001bc01",x"448005bc01",x"448003bc01",x"45000f7c01",x"450000fc01",x"458009fc01",x"458019fc01",x"460027fc01",x"460017fc01",x"46805ffc01",x"46803ffc01",x"3000000000",x"3000000000",x"46807ffc01",x"738001fc00",x"3000000000",
		x"438001f402",x"4380000c02",x"4380010c02",x"440000ec02",x"440002ec02",x"4480033c02",x"4480073c02",x"45800efc02",x"45801efc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458001fc02",x"7280002c00",x"3000000000",
		x"4380008c02",x"4380018c02",x"4380004c02",x"440001ec02",x"440003ec02",x"448000bc02",x"448004bc02",x"458011fc02",x"458009fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458019fc02",x"7280006c00",x"3000000000",
		x"4380014c02",x"4400001c02",x"4400021c02",x"448002bc02",x"448006bc02",x"4500037c02",x"45000b7c02",x"46000bfc02",x"46002bfc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46001bfc02",x"7300003c00",x"3000000000",
		x"4400011c02",x"4400031c02",x"4400009c02",x"448001bc02",x"448005bc02",x"4500077c02",x"45000f7c02",x"46003bfc02",x"460007fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460027fc02",x"730000bc00",x"3000000000",
		x"4300005402",x"438000cc02",x"438001cc02",x"4400029c02",x"4400019c02",x"448003bc02",x"448007bc02",x"458005fc02",x"458015fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45800dfc02",x"7280001c00",x"3000000000",
		x"4380002c02",x"4380012c02",x"438000ac02",x"4400039c02",x"4400005c02",x"4480007c02",x"4480047c02",x"45801dfc02",x"458003fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458013fc02",x"7280005c00",x"3000000000",
		x"4400025c02",x"4400015c02",x"4400035c02",x"4480027c02",x"4480067c02",x"450000fc02",x"450008fc02",x"460017fc02",x"460037fc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46000ffc02",x"7300007c00",x"3000000000",
		x"440000dc02",x"440002dc02",x"440001dc02",x"4480017c02",x"4480057c02",x"450004fc02",x"45000cfc02",x"46002ffc02",x"46001ffc02",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46003ffc02",x"730000fc00",x"3000000000",
		x"4280006403",x"c000000077",x"c000000078",x"4380010c03",x"4380008c03",x"4480063c03",x"4480013c03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480053c03",x"7200002c00",x"3000000000",
		x"430000d403",x"c000000079",x"4380018c03",x"440000ec03",x"440002ec03",x"45000b7c03",x"4500077c03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458006fc03",x"7300005c00",x"3000000000",
		x"4300003403",x"c00000007a",x"4380004c03",x"440001ec03",x"440003ec03",x"45000f7c03",x"450000fc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458016fc03",x"730000dc00",x"3000000000",
		x"4380014c03",x"4400001c03",x"4400021c03",x"4480033c03",x"4480073c03",x"45800efc03",x"45801efc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46002bfc03",x"7380013c00",x"3000000000",
		x"438000cc03",x"4400011c03",x"4400031c03",x"448000bc03",x"448004bc03",x"458001fc03",x"458011fc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46001bfc03",x"738000bc00",x"3000000000",
		x"438001cc03",x"4400009c03",x"4400029c03",x"448002bc03",x"448006bc03",x"458009fc03",x"458019fc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46003bfc03",x"738001bc00",x"3000000000",
		x"4380002c03",x"4400019c03",x"4400039c03",x"448001bc03",x"448005bc03",x"458005fc03",x"458015fc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460007fc03",x"7380007c00",x"3000000000",
		x"4200001404",x"c00000007b",x"4280003404",x"438000cc04",x"438001cc04",x"448007bc04",x"4500057c04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45000d7c04",x"7200000c00",x"3000000000",
		x"c00000007c",x"c00000007d",x"c00000007e",x"4400039c04",x"4400005c04",x"4500037c04",x"45000b7c04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458005fc04",x"7200002c00",x"3000000000",
		x"4280007404",x"c00000007f",x"c000000080",x"4400025c04",x"4400015c04",x"4500077c04",x"458015fc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45800dfc04",x"7280001c00",x"3000000000",
		x"4380002c04",x"4400035c04",x"440000dc04",x"4480007c04",x"45000f7c04",x"46001dfc04",x"46003dfc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468017fc04",x"7300005c00",x"3000000000",
		x"4380012c04",x"440002dc04",x"440001dc04",x"450000fc04",x"450008fc04",x"460003fc04",x"468057fc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468037fc04",x"7380007c00",x"3000000000",
		x"c000000081",x"c000000082",x"c000000083",x"440001ec05",x"448006dc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4500067c05",x"7180001400",x"3000000000",
		x"c000000084",x"c000000085",x"c000000086",x"45000e7c05",x"4500017c05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458002fc05",x"7280000c00",x"3000000000",
		x"c000000087",x"c000000088",x"438000ec05",x"4500097c05",x"4500057c05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460009fc05",x"7280004c00",x"3000000000",
		x"448001dc05",x"45000d7c05",x"4500037c05",x"46803bfc05",x"46807bfc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47002ffc05",x"740000fc00",x"3000000000",
		x"c000000089",x"c00000008a",x"4200001806",x"4400015c06",x"4400035c06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"450000fc06",x"7180000400",x"3000000000",
		x"4200003806",x"c00000008b",x"4300003406",x"450008fc06",x"450004fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46000dfc06",x"7280002c00",x"3000000000",
		x"c00000008c",x"4380006c06",x"4380016c06",x"45800efc06",x"46002dfc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468037fc06",x"7300001c00",x"3000000000",
		x"4200000406",x"c00000008d",x"430000b406",x"45000cfc06",x"450002fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46001dfc06",x"7280006c00",x"3000000000",
		x"c00000008e",x"430000ac07",x"4300006c07",x"460013fc07",x"460033fc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47004ffc07",x"7280002c00",x"3000000000",
		x"4200001407",x"430000ec07",x"c00000008f",x"46000bfc07",x"46002bfc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700cffc07",x"7280006c00",x"3000000000",
		x"c000000090",x"4300001c07",x"4300009c07",x"46001bfc07",x"46003bfc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47002ffc07",x"7280001c00",x"3000000000",
		x"4300005c07",x"440001bc07",x"c000000091",x"4700affc07",x"47006ffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48027ffc07",x"7380007c00",x"3000000000",
		x"c000000092",x"4200003008",x"4200000808",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"450000fc08",x"7180001800",x"3000000000",
		x"4200002808",x"438000ec08",x"438001ec08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46800ffc08",x"7300005c00",x"3000000000",
		x"4200001808",x"4380001c08",x"4380011c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460017fc08",x"730000dc00",x"3000000000",
		x"4380009c08",x"450008fc08",x"450004fc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780bffc08",x"748001fc00",x"3000000000",
		x"4200003808",x"4380019c08",x"4380005c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46804ffc08",x"7380003c00",x"3000000000",
		x"4380015c08",x"45000cfc08",x"450002fc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801fffc08",x"750007fc00",x"3000000000",
		x"c000000093",x"c000000094",x"c000000095",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458013fc09",x"7180000800",x"3000000000",
		x"c000000096",x"4400005c09",x"448003dc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47801ffc09",x"7380001c00",x"3000000000",
		x"c000000097",x"c000000098",x"428000240a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46800ffc0a",x"7180000800",x"3000000000",
		x"c000000099",x"448004bc0a",x"45000ebc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48847ffc0a",x"7400023c00",x"3000000000",
		x"c00000009a",x"448002bc0a",x"450001bc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48827ffc0a",x"7400013c00",x"3000000000",
		x"c00000009b",x"c00000009c",x"430000440b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47006ffc0b",x"7200001000",x"3000000000",
		x"c00000009d",x"4580097c0b",x"4580197c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4981fffc0b",x"7480007c00",x"3000000000",
		x"430000c40b",x"4580057c0b",x"4580157c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a2dfffc0b",x"75000b7c00",x"3000000000",
		x"430000240b",x"45800d7c0b",x"45801d7c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a1dfffc0b",x"7500077c00",x"3000000000",
		x"c00000009e",x"430000c40c",x"c00000009f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780effc0c",x"7200001000",x"3000000000",
		x"c0000000a0",x"460003fc0c",x"468027fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a07fffc0c",x"748000fc00",x"3000000000",
		x"c0000000a1",x"438001840d",x"438000440d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47808ffc0d",x"7280002000",x"3000000000",
		x"438001440d",x"460017fc0d",x"460037fc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490ffffc0d",x"740003fc00",x"3000000000",
		x"c0000000a2",x"440000840e",x"440002840e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48010ffc0e",x"7300004000",x"3000000000",
		x"c0000000a3",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002040f",x"7400010000",x"3000000000",
		x"4380012c03",x"4400005c03",x"4400025c03",x"448003bc03",x"448007bc03",x"45800dfc03",x"45801dfc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460027fc03",x"7380017c00",x"3000000000",
		x"438000ac03",x"4400015c03",x"4400035c03",x"4480007c03",x"4480047c03",x"458003fc03",x"458013fc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460017fc03",x"738000fc00",x"3000000000",
		x"440000dc03",x"4480027c03",x"4480067c03",x"450008fc03",x"450004fc03",x"460037fc03",x"46000ffc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46803ffc03",x"740001fc00",x"3000000000",
		x"440002dc03",x"4480017c03",x"4480057c03",x"45000cfc03",x"450002fc03",x"46002ffc03",x"46001ffc03",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46807ffc03",x"740003fc00",x"3000000000",
		x"4300000c04",x"438000ac04",x"438001ac04",x"4480047c04",x"4480027c04",x"460023fc04",x"460013fc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460033fc04",x"730000dc00",x"3000000000",
		x"4300008c04",x"4380006c04",x"4380016c04",x"4480067c04",x"4480017c04",x"46000bfc04",x"46002bfc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46001bfc04",x"7300003c00",x"3000000000",
		x"438000ec04",x"440003dc04",x"4400003c04",x"450004fc04",x"45000cfc04",x"46003bfc04",x"468077fc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46800ffc04",x"730000bc00",x"3000000000",
		x"438001ec04",x"4400023c04",x"4400013c04",x"450002fc04",x"45000afc04",x"460007fc04",x"46804ffc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46802ffc04",x"7380017c00",x"3000000000",
		x"4380001c04",x"4400033c04",x"440000bc04",x"450006fc04",x"45000efc04",x"460027fc04",x"46806ffc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46801ffc04",x"738000fc00",x"3000000000",
		x"4380011c04",x"440002bc04",x"440001bc04",x"450001fc04",x"450009fc04",x"46805ffc04",x"46803ffc04",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46807ffc04",x"738001fc00",x"3000000000",
		x"4280002c05",x"c0000000a4",x"c0000000a5",x"448005dc05",x"45000b7c05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458012fc05",x"7280002c00",x"3000000000",
		x"c0000000a6",x"440003ec05",x"4400001c05",x"45800afc05",x"45801afc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468007fc05",x"7300006c00",x"3000000000",
		x"c0000000a7",x"4400021c05",x"4400011c05",x"458006fc05",x"458016fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468047fc05",x"730000ec00",x"3000000000",
		x"c0000000a8",x"4400031c05",x"4400009c05",x"45800efc05",x"45801efc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468027fc05",x"7300001c00",x"3000000000",
		x"4400029c05",x"448003dc05",x"448007dc05",x"460029fc05",x"460019fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700affc05",x"738000dc00",x"3000000000",
		x"4400019c05",x"4480003c05",x"4480043c05",x"460039fc05",x"460005fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47006ffc05",x"738001dc00",x"3000000000",
		x"c0000000a9",x"4400039c05",x"4400005c05",x"458001fc05",x"458011fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468067fc05",x"7300009c00",x"3000000000",
		x"4400025c05",x"4480023c05",x"4480063c05",x"460025fc05",x"460015fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700effc05",x"7380003c00",x"3000000000",
		x"4180000806",x"c0000000aa",x"c0000000ab",x"4480017c06",x"4480057c06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45801efc06",x"7200000c00",x"3000000000",
		x"c0000000ac",x"4300007406",x"430000f406",x"45000afc06",x"458001fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"468077fc06",x"7300009c00",x"3000000000",
		x"4300000c06",x"440000dc06",x"440002dc06",x"46003dfc06",x"460003fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47005ffc06",x"738000bc00",x"3000000000",
		x"4300008c06",x"440001dc06",x"440003dc06",x"460023fc06",x"460013fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700dffc06",x"738001bc00",x"3000000000",
		x"c0000000ad",x"4400003c06",x"4400023c06",x"460033fc06",x"46000bfc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47003ffc06",x"7380007c00",x"3000000000",
		x"4200003407",x"c0000000ae",x"c0000000af",x"460007fc07",x"460027fc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700effc07",x"7280005c00",x"3000000000",
		x"438000dc07",x"4480027c07",x"4480067c07",x"47809ffc07",x"47819ffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48017ffc07",x"7400017c00",x"3000000000",
		x"4200000c07",x"c0000000b0",x"c0000000b1",x"460017fc07",x"460037fc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47001ffc07",x"7280003c00",x"3000000000",
		x"4480017c07",x"45801dfc07",x"458003fc07",x"48037ffc07",x"4886fffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490ffffc07",x"748007fc00",x"3000000000",
		x"c0000000b2",x"4200000408",x"c0000000b3",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45000afc08",x"7180000400",x"3000000000",
		x"c0000000b4",x"c0000000b5",x"c0000000b6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45800bfc09",x"7180001800",x"3000000000",
		x"c0000000b7",x"4400025c09",x"4400015c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47811ffc09",x"7380011c00",x"3000000000",
		x"c0000000b8",x"4400035c09",x"448007dc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47809ffc09",x"7380009c00",x"3000000000",
		x"c0000000b9",x"440000dc09",x"4480003c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47819ffc09",x"7380019c00",x"3000000000",
		x"c0000000ba",x"428000640a",x"428000140a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46804ffc0a",x"7180001800",x"3000000000",
		x"428000540a",x"450009bc0a",x"450005bc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48867ffc0a",x"7400033c00",x"3000000000",
		x"428000340a",x"45000dbc0a",x"450003bc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48817ffc0a",x"740000bc00",x"3000000000",
		x"428000740a",x"45000bbc0a",x"450007bc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48857ffc0a",x"740002bc00",x"3000000000",
		x"c0000000bb",x"c0000000bc",x"430000a40b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700effc0b",x"7200003000",x"3000000000",
		x"c0000000bd",x"4580037c0b",x"4580137c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4991fffc0b",x"7480047c00",x"3000000000",
		x"c0000000be",x"45800b7c0b",x"45801b7c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4989fffc0b",x"7480027c00",x"3000000000",
		x"c0000000bf",x"430000240c",x"c0000000c0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781effc0c",x"7200003000",x"3000000000",
		x"c0000000c1",x"460023fc0c",x"468067fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a27fffc0c",x"748004fc00",x"3000000000",
		x"c0000000c2",x"460013fc0c",x"468017fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a17fffc0c",x"748002fc00",x"3000000000",
		x"c0000000c3",x"438000c40d",x"438001c40d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47818ffc0d",x"7280006000",x"3000000000",
		x"c0000000c4",x"440001840e",x"440003840e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48030ffc0e",x"730000c000",x"3000000000",
		x"c0000000c5",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006040f",x"7400030000",x"3000000000",
		x"c0000000c6",x"4480013c05",x"4480053c05",x"460035fc05",x"46000dfc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47001ffc05",x"7380013c00",x"3000000000",
		x"4400015c05",x"4480033c05",x"4480073c05",x"46002dfc05",x"46001dfc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47009ffc05",x"738000bc00",x"3000000000",
		x"c0000000c7",x"448000bc05",x"448004bc05",x"46003dfc05",x"460003fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47005ffc05",x"738001bc00",x"3000000000",
		x"4400035c05",x"448002bc05",x"448006bc05",x"460023fc05",x"460013fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700dffc05",x"7380007c00",x"3000000000",
		x"c0000000c8",x"448001bc05",x"448005bc05",x"460033fc05",x"46000bfc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47003ffc05",x"7300005c00",x"3000000000",
		x"440000dc05",x"448003bc05",x"448007bc05",x"46002bfc05",x"46001bfc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700bffc05",x"7380017c00",x"3000000000",
		x"c0000000c9",x"438000ec06",x"438001ec06",x"458011fc06",x"458009fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46800ffc06",x"7300005c00",x"3000000000",
		x"c0000000ca",x"4380001c06",x"4380011c06",x"458019fc06",x"46002bfc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46804ffc06",x"730000dc00",x"3000000000",
		x"4280005406",x"4380009c06",x"4380019c06",x"458005fc06",x"458015fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46802ffc06",x"7300003c00",x"3000000000",
		x"4380005c06",x"4480037c06",x"4480077c06",x"46806ffc06",x"46801ffc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781fffc06",x"740003fc00",x"3000000000",
		x"438001dc07",x"4480057c07",x"4480037c07",x"47805ffc07",x"47815ffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4881fffc07",x"7400037c00",x"3000000000",
		x"4380003c07",x"4480077c07",x"45000efc07",x"4780dffc07",x"4781dffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4885fffc07",x"740000fc00",x"3000000000",
		x"4380013c07",x"448000fc07",x"448004fc07",x"47803ffc07",x"47813ffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800fffc07",x"740002fc00",x"3000000000",
		x"438000bc07",x"448002fc07",x"450001fc07",x"4780bffc07",x"4781bffc07",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883fffc07",x"740001fc00",x"3000000000",
		x"c0000000cb",x"c0000000cc",x"c0000000cd",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"450006fc08",x"7200001400",x"3000000000",
		x"c0000000ce",x"c0000000cf",x"440001dc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46802ffc08",x"7380013c00",x"3000000000",
		x"c0000000d0",x"c0000000d1",x"4280003809",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45801bfc09",x"7200000400",x"3000000000",
		x"c0000000d2",x"440002dc09",x"4480043c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47805ffc09",x"7380005c00",x"3000000000",
		x"4280007809",x"4480023c09",x"4480063c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800bffc09",x"7400013c00",x"3000000000",
		x"c0000000d3",x"440001dc09",x"4480013c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47815ffc09",x"7380015c00",x"3000000000",
		x"4280000409",x"4480053c09",x"4480033c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802bffc09",x"7400033c00",x"3000000000",
		x"4280004409",x"4480073c09",x"448000bc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780dffc09",x"740000bc00",x"3000000000",
		x"c0000000d4",x"4280000c0a",x"c0000000d5",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46802ffc0a",x"7180000400",x"3000000000",
		x"c0000000d6",x"c0000000d7",x"430000640b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47001ffc0b",x"7200000800",x"3000000000",
		x"c0000000d8",x"4580077c0b",x"4580177c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4999fffc0b",x"7480067c00",x"3000000000",
		x"c0000000d9",x"45800f7c0b",x"45801f7c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4985fffc0b",x"7480017c00",x"3000000000",
		x"c0000000da",x"458000fc0b",x"458010fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4995fffc0b",x"7480057c00",x"3000000000",
		x"c0000000db",x"430000a40c",x"438000540c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47801ffc0c",x"7200000800",x"3000000000",
		x"438001540c",x"460033fc0c",x"468057fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a37fffc0c",x"750007fc00",x"3000000000",
		x"438000d40c",x"46000bfc0c",x"468037fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4abffffc0c",x"75000ffc00",x"3000000000",
		x"438001d40c",x"46002bfc0c",x"468077fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4afffffc0c",x"748006fc00",x"3000000000",
		x"c0000000dc",x"438000240d",x"438001240d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47804ffc0d",x"7280001000",x"3000000000",
		x"c0000000dd",x"440000440e",x"440002440e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48008ffc0e",x"7300002000",x"3000000000",
		x"c0000000de",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001040f",x"7400008000",x"3000000000",
		x"4480007c05",x"4500077c05",x"45000f7c05",x"468017fc05",x"468057fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47007ffc05",x"740002fc00",x"3000000000",
		x"4480047c05",x"450000fc05",x"450008fc05",x"468037fc05",x"468077fc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780fffc05",x"740001fc00",x"3000000000",
		x"4480027c05",x"450004fc05",x"45000cfc05",x"46800ffc05",x"46804ffc05",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781fffc05",x"740003fc00",x"3000000000",
		x"4300004c06",x"4400013c06",x"4400033c06",x"46001bfc06",x"46003bfc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700bffc06",x"7380017c00",x"3000000000",
		x"430000cc06",x"440000bc06",x"440002bc06",x"460007fc06",x"460027fc06",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47007ffc06",x"738000fc00",x"3000000000",
		x"c0000000df",x"4280002408",x"4280006408",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45800dfc08",x"7200003400",x"3000000000",
		x"4280001408",x"440003dc08",x"4400003c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46806ffc08",x"738000bc00",x"3000000000",
		x"4280005408",x"4400023c08",x"4400013c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47001ffc08",x"7400007c00",x"3000000000",
		x"4280003408",x"4400033c08",x"440000bc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47009ffc08",x"738001bc00",x"3000000000",
		x"440002bc08",x"45801dfc08",x"458003fc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803fffc08",x"75000ffc00",x"3000000000",
		x"c0000000e0",x"4280002409",x"4280006409",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460007fc09",x"7200002400",x"3000000000",
		x"4280001409",x"448004bc09",x"448002bc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781dffc09",x"738000dc00",x"3000000000",
		x"4280005409",x"448006bc09",x"448001bc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47803ffc09",x"738001dc00",x"3000000000",
		x"4280003409",x"448005bc09",x"448003bc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47813ffc09",x"7380003c00",x"3000000000",
		x"c0000000e1",x"4280004c0a",x"c0000000e2",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46806ffc0a",x"7180001400",x"3000000000",
		x"c0000000e3",x"45000fbc0a",x"4500007c0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48837ffc0a",x"740001bc00",x"3000000000",
		x"c0000000e4",x"c0000000e5",x"430000e40b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47009ffc0b",x"7200002800",x"3000000000",
		x"c0000000e6",x"458008fc0b",x"458018fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a3dfffc0b",x"75000f7c00",x"3000000000",
		x"c0000000e7",x"458004fc0b",x"458014fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a03fffc0b",x"750000fc00",x"3000000000",
		x"c0000000e8",x"45800cfc0b",x"45801cfc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a23fffc0b",x"750008fc00",x"3000000000",
		x"c0000000e9",x"458002fc0b",x"458012fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a13fffc0b",x"750004fc00",x"3000000000",
		x"c0000000ea",x"430000640c",x"438000340c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47811ffc0c",x"7280002800",x"3000000000",
		x"c0000000eb",x"438000a40d",x"438001a40d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47814ffc0d",x"7280005000",x"3000000000",
		x"c0000000ec",x"440001440e",x"440003440e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48028ffc0e",x"730000a000",x"3000000000",
		x"c0000000ed",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005040f",x"7400028000",x"3000000000",
		x"c0000000ee",x"4280007408",x"c0000000ef",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"458013fc08",x"7280000c00",x"3000000000",
		x"c0000000f0",x"4280007409",x"c0000000f1",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460027fc09",x"7200001400",x"3000000000",
		x"c0000000f2",x"4280002c0a",x"c0000000f3",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46801ffc0a",x"7200000c00",x"3000000000",
		x"c0000000f4",x"4500087c0a",x"4500047c0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"49077ffc0a",x"748003bc00",x"3000000000",
		x"c0000000f5",x"45000c7c0a",x"4500027c0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490f7ffc0a",x"748007bc00",x"3000000000",
		x"c0000000f6",x"c0000000f7",x"430000140b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47005ffc0b",x"7200001800",x"3000000000",
		x"c0000000f8",x"45800afc0b",x"45801afc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a33fffc0b",x"75000cfc00",x"3000000000",
		x"430000940b",x"458006fc0b",x"458016fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a0bfffc0b",x"750002fc00",x"3000000000",
		x"430000540b",x"45800efc0b",x"45801efc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a2bfffc0b",x"75000afc00",x"3000000000",
		x"430000d40b",x"458001fc0b",x"458011fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a1bfffc0b",x"750006fc00",x"3000000000",
		x"c0000000f9",x"458009fc0b",x"458019fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a3bfffc0b",x"75000efc00",x"3000000000",
		x"c0000000fa",x"430000e40c",x"438001340c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47809ffc0c",x"7280006800",x"3000000000",
		x"c0000000fb",x"438000640d",x"438001640d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780cffc0d",x"7280003000",x"3000000000",
		x"c0000000fc",x"440000c40e",x"440002c40e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48018ffc0e",x"7300006000",x"3000000000",
		x"c0000000fd",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003040f",x"7400018000",x"3000000000",
		x"c0000000fe",x"c0000000ff",x"c000000100",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45800bfc08",x"7280004c00",x"3000000000",
		x"c000000101",x"448003bc08",x"448007bc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47005ffc08",x"7400027c00",x"3000000000",
		x"c000000102",x"4280000c09",x"c000000103",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460017fc09",x"7200003400",x"3000000000",
		x"c000000104",x"448007bc09",x"4500097c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801bffc09",x"740002bc00",x"3000000000",
		x"c000000105",x"c000000106",x"c000000107",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46805ffc0a",x"7200002c00",x"3000000000",
		x"c000000108",x"45000a7c0a",x"458001fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4900fffc0a",x"7480007c00",x"3000000000",
		x"c000000109",x"4500067c0a",x"458011fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4908fffc0a",x"7480047c00",x"3000000000",
		x"c00000010a",x"45000e7c0a",x"458009fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4904fffc0a",x"7480027c00",x"3000000000",
		x"c00000010b",x"430000340b",x"430000b40b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780dffc0b",x"7200003800",x"3000000000",
		x"430000740b",x"458005fc0b",x"458015fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a07fffc0b",x"750001fc00",x"3000000000",
		x"430000f40b",x"45800dfc0b",x"45801dfc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a27fffc0b",x"750009fc00",x"3000000000",
		x"4300000c0b",x"458003fc0b",x"460013fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a17fffc0b",x"750005fc00",x"3000000000",
		x"c00000010c",x"430000140c",x"438000b40c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47819ffc0c",x"7280001800",x"3000000000",
		x"c00000010d",x"438000e40d",x"438001e40d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781cffc0d",x"7280007000",x"3000000000",
		x"c00000010e",x"440001c40e",x"440003c40e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48038ffc0e",x"730000e000",x"3000000000",
		x"c00000010f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007040f",x"7400038000",x"3000000000",
		x"c000000110",x"4300000c08",x"4300008c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"45801bfc08",x"7280002c00",x"3000000000",
		x"c000000111",x"4480007c08",x"4480047c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4700dffc08",x"7400017c00",x"3000000000",
		x"4300004c08",x"4480027c08",x"4480067c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781bffc08",x"7400037c00",x"3000000000",
		x"430000cc08",x"4480017c08",x"4480057c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47003ffc08",x"740000fc00",x"3000000000",
		x"c000000112",x"c000000113",x"c000000114",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460037fc09",x"7200000c00",x"3000000000",
		x"c000000115",x"4480007c09",x"4500057c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803bffc09",x"740001bc00",x"3000000000",
		x"c000000116",x"4480047c09",x"45000d7c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48007ffc09",x"740003bc00",x"3000000000",
		x"408000000a",x"c000000117",x"c000000118",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46803ffc0a",x"7200001c00",x"3000000000",
		x"c000000119",x"4500017c0a",x"4500097c0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490cfffc0a",x"7480067c00",x"3000000000",
		x"c00000011a",x"4500057c0a",x"458019fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4902fffc0a",x"7480017c00",x"3000000000",
		x"4300006c0a",x"45000d7c0a",x"458005fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490afffc0a",x"7480057c00",x"3000000000",
		x"430000ec0a",x"4500037c0a",x"458015fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4906fffc0a",x"7480037c00",x"3000000000",
		x"4300001c0a",x"45000b7c0a",x"45800dfc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490efffc0a",x"7480077c00",x"3000000000",
		x"c00000011b",x"4300008c0b",x"4300004c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781dffc0b",x"7200000400",x"3000000000",
		x"c00000011c",x"430000940c",x"438001b40c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47805ffc0c",x"7280005800",x"3000000000",
		x"c00000011d",x"438000140d",x"438001140d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47802ffc0d",x"7280000800",x"3000000000",
		x"c00000011e",x"440000240e",x"440002240e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48004ffc0e",x"7300001000",x"3000000000",
		x"c00000011f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000840f",x"7400004000",x"3000000000",
		x"4180000008",x"4300002c08",x"c000000120",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"460037fc08",x"7280006c00",x"3000000000",
		x"430000ac08",x"4480037c08",x"4480077c08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47807ffc08",x"740002fc00",x"3000000000",
		x"c000000121",x"c000000122",x"4300004c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46000ffc09",x"7280002c00",x"3000000000",
		x"c000000123",x"4480027c09",x"4500037c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48027ffc09",x"7400007c00",x"3000000000",
		x"430000cc09",x"45000b7c09",x"4500077c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4881fffc09",x"7400027c00",x"3000000000",
		x"4300002c09",x"45000f7c09",x"450000fc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48017ffc09",x"7400017c00",x"3000000000",
		x"430000ac09",x"450008fc09",x"450004fc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48037ffc09",x"7400037c00",x"3000000000",
		x"c000000124",x"4500077c0a",x"45000f7c0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4901fffc0a",x"748000fc00",x"3000000000",
		x"4300009c0a",x"450000fc0a",x"45801dfc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4909fffc0a",x"748004fc00",x"3000000000",
		x"c000000125",x"450008fc0a",x"450004fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4905fffc0a",x"748002fc00",x"3000000000",
		x"4300005c0a",x"45000cfc0a",x"458003fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490dfffc0a",x"748006fc00",x"3000000000",
		x"c000000126",x"430000cc0b",x"4300002c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47803ffc0b",x"7200002400",x"3000000000",
		x"c000000127",x"c000000128",x"438000740c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47815ffc0c",x"7280003800",x"3000000000",
		x"c000000129",x"438000940d",x"4400004c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47812ffc0d",x"7280004800",x"3000000000",
		x"c00000012a",x"440001240e",x"440003240e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48024ffc0e",x"7300009000",x"3000000000",
		x"c00000012b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004840f",x"7400024000",x"3000000000",
		x"c00000012c",x"45000efc08",x"450001fc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47817ffc08",x"748005fc00",x"3000000000",
		x"4100000009",x"c00000012d",x"4300006c09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"46002ffc09",x"7280006c00",x"3000000000",
		x"c00000012e",x"45000cfc09",x"450002fc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800fffc09",x"740000fc00",x"3000000000",
		x"c00000012f",x"4480067c09",x"45000afc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802fffc09",x"740002fc00",x"3000000000",
		x"c000000130",x"450002fc0a",x"458013fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4903fffc0a",x"748001fc00",x"3000000000",
		x"c000000131",x"45000afc0a",x"45800bfc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490bfffc0a",x"748005fc00",x"3000000000",
		x"c000000132",x"430000ac0b",x"4300006c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47813ffc0b",x"7200001400",x"3000000000",
		x"c000000133",x"c000000134",x"438001740c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780dffc0c",x"7280007800",x"3000000000",
		x"c000000135",x"46001bfc0c",x"46800ffc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a0ffffc0c",x"748001fc00",x"3000000000",
		x"c000000136",x"438001940d",x"4400024c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780affc0d",x"7280002800",x"3000000000",
		x"c000000137",x"440000a40e",x"440002a40e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48014ffc0e",x"7300005000",x"3000000000",
		x"c000000138",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002840f",x"7400014000",x"3000000000",
		x"438000dc08",x"450009fc08",x"450005fc08",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780fffc08",x"748003fc00",x"3000000000",
		x"430000ec09",x"450006fc09",x"45000efc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4885fffc09",x"748003fc00",x"3000000000",
		x"4300001c09",x"450001fc09",x"450009fc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883fffc09",x"748007fc00",x"3000000000",
		x"4300009c09",x"450005fc09",x"45000dfc09",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4887fffc09",x"740001fc00",x"3000000000",
		x"430000dc0a",x"450006fc0a",x"45801bfc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4907fffc0a",x"748003fc00",x"3000000000",
		x"4300003c0a",x"45000efc0a",x"458007fc0a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"490ffffc0a",x"748007fc00",x"3000000000",
		x"c000000139",x"430000ec0b",x"c00000013a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780bffc0b",x"7200003400",x"3000000000",
		x"c00000013b",x"438000f40c",x"438001f40c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781dffc0c",x"7280000400",x"3000000000",
		x"4380000c0c",x"46003bfc0c",x"46804ffc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a2ffffc0c",x"748005fc00",x"3000000000",
		x"4380010c0c",x"460007fc0c",x"46802ffc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a1ffffc0c",x"748003fc00",x"3000000000",
		x"c00000013c",x"438000540d",x"4400014c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781affc0d",x"7280006800",x"3000000000",
		x"c00000013d",x"440001a40e",x"440003a40e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48034ffc0e",x"730000d000",x"3000000000",
		x"c00000013e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006840f",x"7400034000",x"3000000000",
		x"c00000013f",x"4300001c0b",x"c000000140",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781bffc0b",x"7200000c00",x"3000000000",
		x"c000000141",x"460033fc0b",x"46000bfc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a37fffc0b",x"75000dfc00",x"3000000000",
		x"c000000142",x"4380008c0c",x"4380018c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47803ffc0c",x"7280004400",x"3000000000",
		x"c000000143",x"438001540d",x"4400034c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47806ffc0d",x"7280001800",x"3000000000",
		x"c000000144",x"440000640e",x"440002640e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800cffc0e",x"7300003000",x"3000000000",
		x"c000000145",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001840f",x"740000c000",x"3000000000",
		x"c000000146",x"4300009c0b",x"c000000147",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47807ffc0b",x"7200002c00",x"3000000000",
		x"4380003c0b",x"46002bfc0b",x"46001bfc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a0ffffc0b",x"750003fc00",x"3000000000",
		x"c000000148",x"46003bfc0b",x"460007fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a2ffffc0b",x"75000bfc00",x"3000000000",
		x"c000000149",x"4380004c0c",x"4380014c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48013ffc0c",x"7280002400",x"3000000000",
		x"c00000014a",x"438000d40d",x"440000cc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47816ffc0d",x"7280005800",x"3000000000",
		x"c00000014b",x"440001640e",x"440003640e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802cffc0e",x"730000b000",x"3000000000",
		x"c00000014c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005840f",x"740002c000",x"3000000000",
		x"c00000014d",x"4300005c0b",x"4380013c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47817ffc0b",x"7200001c00",x"3000000000",
		x"438000bc0b",x"460027fc0b",x"460017fc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a1ffffc0b",x"750007fc00",x"3000000000",
		x"438001bc0b",x"460037fc0b",x"46000ffc0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4a3ffffc0b",x"75000ffc00",x"3000000000",
		x"c00000014e",x"438000cc0c",x"438001cc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48033ffc0c",x"7280006400",x"3000000000",
		x"c00000014f",x"438001d40d",x"440002cc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780effc0d",x"7280003800",x"3000000000",
		x"c000000150",x"440000e40e",x"440002e40e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801cffc0e",x"7300007000",x"3000000000",
		x"c000000151",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003840f",x"740001c000",x"3000000000",
		x"408000000b",x"430000dc0b",x"4380007c0b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4780fffc0b",x"7280003c00",x"3000000000",
		x"c000000152",x"4380002c0c",x"4380012c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800bffc0c",x"7280001400",x"3000000000",
		x"c000000153",x"438000340d",x"440001cc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4781effc0d",x"7280007800",x"3000000000",
		x"c000000154",x"440001e40e",x"440003e40e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803cffc0e",x"730000f000",x"3000000000",
		x"c000000155",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007840f",x"740003c000",x"3000000000",
		x"c000000156",x"438000ac0c",x"438001ac0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802bffc0c",x"7280005400",x"3000000000",
		x"c000000157",x"438001340d",x"440003cc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47801ffc0d",x"7280000400",x"3000000000",
		x"c000000158",x"440000140e",x"440002140e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48002ffc0e",x"7300000800",x"3000000000",
		x"c000000159",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000440f",x"7400002000",x"3000000000",
		x"c00000015a",x"4380006c0c",x"4380016c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801bffc0c",x"7280003400",x"3000000000",
		x"c00000015b",x"438000b40d",x"4400002c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"47811ffc0d",x"7280004400",x"3000000000",
		x"c00000015c",x"440001140e",x"440003140e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48022ffc0e",x"7300008800",x"3000000000",
		x"c00000015d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004440f",x"7400022000",x"3000000000",
		x"c00000015e",x"438000ec0c",x"438001ec0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803bffc0c",x"7280007400",x"3000000000",
		x"c00000015f",x"438001b40d",x"4400022c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48009ffc0d",x"7300002400",x"3000000000",
		x"c000000160",x"440000940e",x"440002940e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48012ffc0e",x"7300004800",x"3000000000",
		x"c000000161",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002440f",x"7400012000",x"3000000000",
		x"c000000162",x"4380001c0c",x"4380011c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48007ffc0c",x"7280000c00",x"3000000000",
		x"c000000163",x"438000740d",x"4400012c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48029ffc0d",x"730000a400",x"3000000000",
		x"c000000164",x"440001940e",x"440003940e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48032ffc0e",x"730000c800",x"3000000000",
		x"c000000165",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006440f",x"7400032000",x"3000000000",
		x"c000000166",x"4380009c0c",x"4380019c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48027ffc0c",x"7280004c00",x"3000000000",
		x"c000000167",x"438001740d",x"4400032c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48019ffc0d",x"7300006400",x"3000000000",
		x"c000000168",x"440000540e",x"440002540e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800affc0e",x"7300002800",x"3000000000",
		x"c000000169",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001440f",x"740000a000",x"3000000000",
		x"c00000016a",x"4380005c0c",x"4380015c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48017ffc0c",x"7280002c00",x"3000000000",
		x"c00000016b",x"438000f40d",x"440000ac0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48039ffc0d",x"730000e400",x"3000000000",
		x"c00000016c",x"440001540e",x"448001ac0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802affc0e",x"730000a800",x"3000000000",
		x"c00000016d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005440f",x"740002a000",x"3000000000",
		x"c00000016e",x"438000dc0c",x"438001dc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48037ffc0c",x"7280006c00",x"3000000000",
		x"c00000016f",x"438001f40d",x"440002ac0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48005ffc0d",x"7300001400",x"3000000000",
		x"c000000170",x"440003540e",x"448005ac0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801affc0e",x"7300006800",x"3000000000",
		x"c000000171",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003440f",x"740001a000",x"3000000000",
		x"c000000172",x"4380003c0c",x"4380013c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800fffc0c",x"7280001c00",x"3000000000",
		x"c000000173",x"4380000c0d",x"440001ac0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48025ffc0d",x"7300009400",x"3000000000",
		x"c000000174",x"440000d40e",x"448003ac0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803affc0e",x"730000e800",x"3000000000",
		x"c000000175",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007440f",x"740003a000",x"3000000000",
		x"c000000176",x"438000bc0c",x"438001bc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802fffc0c",x"7280005c00",x"3000000000",
		x"c000000177",x"4380010c0d",x"440003ac0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48015ffc0d",x"7300005400",x"3000000000",
		x"c000000178",x"440002d40e",x"448007ac0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48006ffc0e",x"7300001800",x"3000000000",
		x"c000000179",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000c40f",x"7400006000",x"3000000000",
		x"c00000017a",x"4380007c0c",x"4380017c0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801fffc0c",x"7280003c00",x"3000000000",
		x"c00000017b",x"4380008c0d",x"4400006c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48035ffc0d",x"730000d400",x"3000000000",
		x"c00000017c",x"440001d40e",x"4480006c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48026ffc0e",x"7300009800",x"3000000000",
		x"c00000017d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004c40f",x"7400026000",x"3000000000",
		x"408000000c",x"438000fc0c",x"440001fc0c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883fffc0c",x"7300007c00",x"3000000000",
		x"c00000017e",x"4380018c0d",x"4400026c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800dffc0d",x"7300003400",x"3000000000",
		x"c00000017f",x"440003d40e",x"4480046c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48016ffc0e",x"7300005800",x"3000000000",
		x"c000000180",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002c40f",x"7400016000",x"3000000000",
		x"c000000181",x"4400016c0d",x"4400036c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802dffc0d",x"730000b400",x"3000000000",
		x"c000000182",x"440000340e",x"4480026c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48036ffc0e",x"730000d800",x"3000000000",
		x"c000000183",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006c40f",x"7400036000",x"3000000000",
		x"c000000184",x"440000ec0d",x"440002ec0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801dffc0d",x"7300007400",x"3000000000",
		x"c000000185",x"440002340e",x"4480066c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800effc0e",x"7300003800",x"3000000000",
		x"c000000186",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001c40f",x"740000e000",x"3000000000",
		x"c000000187",x"440001ec0d",x"440003ec0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803dffc0d",x"730000f400",x"3000000000",
		x"c000000188",x"440001340e",x"4480016c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802effc0e",x"730000b800",x"3000000000",
		x"c000000189",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005c40f",x"740002e000",x"3000000000",
		x"c00000018a",x"4400001c0d",x"4400021c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48003ffc0d",x"7300000c00",x"3000000000",
		x"c00000018b",x"440003340e",x"4480056c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801effc0e",x"7300007800",x"3000000000",
		x"c00000018c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003c40f",x"740001e000",x"3000000000",
		x"c00000018d",x"4400011c0d",x"4400031c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48023ffc0d",x"7300008c00",x"3000000000",
		x"c00000018e",x"440000b40e",x"4480036c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803effc0e",x"730000f800",x"3000000000",
		x"c00000018f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007c40f",x"740003e000",x"3000000000",
		x"c000000190",x"4400009c0d",x"4400029c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48013ffc0d",x"7300004c00",x"3000000000",
		x"c000000191",x"440002b40e",x"4480076c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48001ffc0e",x"7300000400",x"3000000000",
		x"c000000192",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000240f",x"7400001000",x"3000000000",
		x"c000000193",x"4400019c0d",x"4400039c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48033ffc0d",x"730000cc00",x"3000000000",
		x"c000000194",x"440001b40e",x"448000ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48021ffc0e",x"7300008400",x"3000000000",
		x"c000000195",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004240f",x"7400021000",x"3000000000",
		x"c000000196",x"4400005c0d",x"4400025c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800bffc0d",x"7300002c00",x"3000000000",
		x"c000000197",x"440003b40e",x"448004ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48011ffc0e",x"7300004400",x"3000000000",
		x"c000000198",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002240f",x"7400011000",x"3000000000",
		x"c000000199",x"4400015c0d",x"4400035c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802bffc0d",x"730000ac00",x"3000000000",
		x"c00000019a",x"440000740e",x"448002ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48031ffc0e",x"730000c400",x"3000000000",
		x"c00000019b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006240f",x"7400031000",x"3000000000",
		x"c00000019c",x"440000dc0d",x"440002dc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801bffc0d",x"7300006c00",x"3000000000",
		x"c00000019d",x"440002740e",x"448006ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48009ffc0e",x"7300002400",x"3000000000",
		x"c00000019e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001240f",x"7400009000",x"3000000000",
		x"c00000019f",x"440001dc0d",x"440003dc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4803bffc0d",x"730000ec00",x"3000000000",
		x"c0000001a0",x"440001740e",x"448001ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48029ffc0e",x"730000a400",x"3000000000",
		x"c0000001a1",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005240f",x"7400029000",x"3000000000",
		x"c0000001a2",x"4400003c0d",x"4400023c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48007ffc0d",x"7300001c00",x"3000000000",
		x"c0000001a3",x"440003740e",x"448005ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48019ffc0e",x"7300006400",x"3000000000",
		x"c0000001a4",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003240f",x"7400019000",x"3000000000",
		x"c0000001a5",x"4400013c0d",x"4400033c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48027ffc0d",x"7300009c00",x"3000000000",
		x"c0000001a6",x"440000f40e",x"448003ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48039ffc0e",x"730000e400",x"3000000000",
		x"c0000001a7",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007240f",x"7400039000",x"3000000000",
		x"c0000001a8",x"440000bc0d",x"440002bc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48017ffc0d",x"7300005c00",x"3000000000",
		x"c0000001a9",x"440002f40e",x"448007ec0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48005ffc0e",x"7300001400",x"3000000000",
		x"c0000001aa",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000a40f",x"7400005000",x"3000000000",
		x"c0000001ab",x"440001bc0d",x"440003bc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48037ffc0d",x"730000dc00",x"3000000000",
		x"c0000001ac",x"440001f40e",x"4480001c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48025ffc0e",x"7300009400",x"3000000000",
		x"c0000001ad",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004a40f",x"7400025000",x"3000000000",
		x"c0000001ae",x"4400007c0d",x"4400027c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4800fffc0d",x"7300003c00",x"3000000000",
		x"c0000001af",x"440003f40e",x"4480041c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48015ffc0e",x"7300005400",x"3000000000",
		x"c0000001b0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002a40f",x"7400015000",x"3000000000",
		x"c0000001b1",x"4400017c0d",x"4400037c0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4802fffc0d",x"730000bc00",x"3000000000",
		x"c0000001b2",x"4400000c0e",x"4480021c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48835ffc0e",x"738000d400",x"3000000000",
		x"c0000001b3",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006a40f",x"7400035000",x"3000000000",
		x"c0000001b4",x"440000fc0d",x"440002fc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4801fffc0d",x"7300007c00",x"3000000000",
		x"c0000001b5",x"4400020c0e",x"4480061c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48875ffc0e",x"738001d400",x"3000000000",
		x"c0000001b6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001a40f",x"740000d000",x"3000000000",
		x"408000000d",x"440001fc0d",x"448003fc0d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883fffc0d",x"738000fc00",x"3000000000",
		x"c0000001b7",x"4400010c0e",x"4480011c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4880dffc0e",x"7380003400",x"3000000000",
		x"c0000001b8",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005a40f",x"740002d000",x"3000000000",
		x"c0000001b9",x"4400030c0e",x"4480051c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4884dffc0e",x"7380013400",x"3000000000",
		x"c0000001ba",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003a40f",x"740001d000",x"3000000000",
		x"c0000001bb",x"4400008c0e",x"4480031c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4882dffc0e",x"738000b400",x"3000000000",
		x"c0000001bc",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007a40f",x"740003d000",x"3000000000",
		x"c0000001bd",x"4400028c0e",x"4480071c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4886dffc0e",x"738001b400",x"3000000000",
		x"c0000001be",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000640f",x"7400003000",x"3000000000",
		x"c0000001bf",x"4400018c0e",x"4480009c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4881dffc0e",x"7380007400",x"3000000000",
		x"c0000001c0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004640f",x"7400023000",x"3000000000",
		x"c0000001c1",x"4400038c0e",x"4480049c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4885dffc0e",x"7380017400",x"3000000000",
		x"c0000001c2",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002640f",x"7400013000",x"3000000000",
		x"c0000001c3",x"4400004c0e",x"4480029c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883dffc0e",x"738000f400",x"3000000000",
		x"c0000001c4",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006640f",x"7400033000",x"3000000000",
		x"c0000001c5",x"4400024c0e",x"4480069c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4887dffc0e",x"738001f400",x"3000000000",
		x"c0000001c6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001640f",x"740000b000",x"3000000000",
		x"c0000001c7",x"4400014c0e",x"4480019c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48803ffc0e",x"7380000c00",x"3000000000",
		x"c0000001c8",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005640f",x"740002b000",x"3000000000",
		x"c0000001c9",x"4400034c0e",x"4480059c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48843ffc0e",x"7380010c00",x"3000000000",
		x"c0000001ca",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003640f",x"740001b000",x"3000000000",
		x"c0000001cb",x"440000cc0e",x"4480039c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48823ffc0e",x"7380008c00",x"3000000000",
		x"c0000001cc",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007640f",x"740003b000",x"3000000000",
		x"c0000001cd",x"440002cc0e",x"4480079c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48863ffc0e",x"7380018c00",x"3000000000",
		x"c0000001ce",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000e40f",x"7400007000",x"3000000000",
		x"c0000001cf",x"440001cc0e",x"4480005c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48813ffc0e",x"7380004c00",x"3000000000",
		x"c0000001d0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004e40f",x"7400027000",x"3000000000",
		x"c0000001d1",x"440003cc0e",x"4480045c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48853ffc0e",x"7380014c00",x"3000000000",
		x"c0000001d2",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002e40f",x"7400017000",x"3000000000",
		x"c0000001d3",x"4400002c0e",x"4480025c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48833ffc0e",x"738000cc00",x"3000000000",
		x"c0000001d4",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006e40f",x"7400037000",x"3000000000",
		x"c0000001d5",x"4400022c0e",x"4480065c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48873ffc0e",x"738001cc00",x"3000000000",
		x"c0000001d6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001e40f",x"740000f000",x"3000000000",
		x"c0000001d7",x"4400012c0e",x"4480015c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4880bffc0e",x"7380002c00",x"3000000000",
		x"c0000001d8",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005e40f",x"740002f000",x"3000000000",
		x"c0000001d9",x"4400032c0e",x"4480055c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4884bffc0e",x"7380012c00",x"3000000000",
		x"c0000001da",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003e40f",x"740001f000",x"3000000000",
		x"c0000001db",x"440000ac0e",x"4480035c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4882bffc0e",x"738000ac00",x"3000000000",
		x"c0000001dc",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007e40f",x"740003f000",x"3000000000",
		x"c0000001dd",x"440002ac0e",x"4480075c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4886bffc0e",x"738001ac00",x"3000000000",
		x"c0000001de",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000140f",x"7400000800",x"3000000000",
		x"c0000001df",x"448000dc0e",x"448004dc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4881bffc0e",x"7380006c00",x"3000000000",
		x"c0000001e0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004140f",x"7400020800",x"3000000000",
		x"c0000001e1",x"448002dc0e",x"448006dc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4885bffc0e",x"7380016c00",x"3000000000",
		x"c0000001e2",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002140f",x"7400010800",x"3000000000",
		x"c0000001e3",x"448001dc0e",x"448005dc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883bffc0e",x"738000ec00",x"3000000000",
		x"c0000001e4",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006140f",x"7400030800",x"3000000000",
		x"c0000001e5",x"448003dc0e",x"448007dc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4887bffc0e",x"738001ec00",x"3000000000",
		x"c0000001e6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001140f",x"7400008800",x"3000000000",
		x"c0000001e7",x"4480003c0e",x"4480043c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48807ffc0e",x"7380001c00",x"3000000000",
		x"c0000001e8",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005140f",x"7400028800",x"3000000000",
		x"c0000001e9",x"4480023c0e",x"4480063c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48847ffc0e",x"7380011c00",x"3000000000",
		x"c0000001ea",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003140f",x"7400018800",x"3000000000",
		x"c0000001eb",x"4480013c0e",x"4480053c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48827ffc0e",x"7380009c00",x"3000000000",
		x"c0000001ec",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007140f",x"7400038800",x"3000000000",
		x"c0000001ed",x"4480033c0e",x"4480073c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48867ffc0e",x"7380019c00",x"3000000000",
		x"c0000001ee",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000940f",x"7400004800",x"3000000000",
		x"c0000001ef",x"448000bc0e",x"448004bc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48817ffc0e",x"7380005c00",x"3000000000",
		x"c0000001f0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004940f",x"7400024800",x"3000000000",
		x"c0000001f1",x"448002bc0e",x"448006bc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48857ffc0e",x"7380015c00",x"3000000000",
		x"c0000001f2",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002940f",x"7400014800",x"3000000000",
		x"c0000001f3",x"448001bc0e",x"448005bc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48837ffc0e",x"738000dc00",x"3000000000",
		x"c0000001f4",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006940f",x"7400034800",x"3000000000",
		x"c0000001f5",x"448003bc0e",x"448007bc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"48877ffc0e",x"738001dc00",x"3000000000",
		x"c0000001f6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001940f",x"740000c800",x"3000000000",
		x"c0000001f7",x"4480007c0e",x"4480047c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4880fffc0e",x"7380003c00",x"3000000000",
		x"c0000001f8",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005940f",x"740002c800",x"3000000000",
		x"c0000001f9",x"4480027c0e",x"4480067c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4884fffc0e",x"7380013c00",x"3000000000",
		x"c0000001fa",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003940f",x"740001c800",x"3000000000",
		x"c0000001fb",x"4480017c0e",x"4480057c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4882fffc0e",x"738000bc00",x"3000000000",
		x"c0000001fc",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007940f",x"740003c800",x"3000000000",
		x"c0000001fd",x"4480037c0e",x"4480077c0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4886fffc0e",x"738001bc00",x"3000000000",
		x"c0000001fe",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000540f",x"7400002800",x"3000000000",
		x"c0000001ff",x"448000fc0e",x"448004fc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4881fffc0e",x"7380007c00",x"3000000000",
		x"c000000200",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004540f",x"7400022800",x"3000000000",
		x"c000000201",x"448002fc0e",x"448006fc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4885fffc0e",x"7380017c00",x"3000000000",
		x"c000000202",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002540f",x"7400012800",x"3000000000",
		x"c000000203",x"448001fc0e",x"448005fc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4883fffc0e",x"738000fc00",x"3000000000",
		x"c000000204",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006540f",x"7400032800",x"3000000000",
		x"408000000e",x"448003fc0e",x"450007fc0e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4887fffc0e",x"738001fc00",x"3000000000",
		x"c000000205",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001540f",x"740000a800",x"3000000000",
		x"c000000206",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005540f",x"740002a800",x"3000000000",
		x"c000000207",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003540f",x"740001a800",x"3000000000",
		x"c000000208",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007540f",x"740003a800",x"3000000000",
		x"c000000209",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000d40f",x"7400006800",x"3000000000",
		x"c00000020a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004d40f",x"7400026800",x"3000000000",
		x"c00000020b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002d40f",x"7400016800",x"3000000000",
		x"c00000020c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006d40f",x"7400036800",x"3000000000",
		x"c00000020d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001d40f",x"740000e800",x"3000000000",
		x"c00000020e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005d40f",x"740002e800",x"3000000000",
		x"c00000020f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003d40f",x"740001e800",x"3000000000",
		x"c000000210",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007d40f",x"740003e800",x"3000000000",
		x"c000000211",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000340f",x"7400001800",x"3000000000",
		x"c000000212",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004340f",x"7400021800",x"3000000000",
		x"c000000213",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002340f",x"7400011800",x"3000000000",
		x"c000000214",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006340f",x"7400031800",x"3000000000",
		x"c000000215",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001340f",x"7400009800",x"3000000000",
		x"c000000216",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005340f",x"7400029800",x"3000000000",
		x"c000000217",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003340f",x"7400019800",x"3000000000",
		x"c000000218",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007340f",x"7400039800",x"3000000000",
		x"c000000219",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000b40f",x"7400005800",x"3000000000",
		x"c00000021a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004b40f",x"7400025800",x"3000000000",
		x"c00000021b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002b40f",x"7400015800",x"3000000000",
		x"c00000021c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006b40f",x"7400035800",x"3000000000",
		x"c00000021d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001b40f",x"740000d800",x"3000000000",
		x"c00000021e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005b40f",x"740002d800",x"3000000000",
		x"c00000021f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003b40f",x"740001d800",x"3000000000",
		x"c000000220",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007b40f",x"740003d800",x"3000000000",
		x"c000000221",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000740f",x"7400003800",x"3000000000",
		x"c000000222",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004740f",x"7400023800",x"3000000000",
		x"c000000223",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002740f",x"7400013800",x"3000000000",
		x"c000000224",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006740f",x"7400033800",x"3000000000",
		x"c000000225",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001740f",x"740000b800",x"3000000000",
		x"c000000226",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005740f",x"740002b800",x"3000000000",
		x"c000000227",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003740f",x"740001b800",x"3000000000",
		x"c000000228",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007740f",x"740003b800",x"3000000000",
		x"c000000229",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000f40f",x"7400007800",x"3000000000",
		x"c00000022a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004f40f",x"7400027800",x"3000000000",
		x"c00000022b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002f40f",x"7400017800",x"3000000000",
		x"c00000022c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006f40f",x"7400037800",x"3000000000",
		x"c00000022d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001f40f",x"740000f800",x"3000000000",
		x"c00000022e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005f40f",x"740002f800",x"3000000000",
		x"c00000022f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003f40f",x"740001f800",x"3000000000",
		x"c000000230",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007f40f",x"740003f800",x"3000000000",
		x"c000000231",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480000c0f",x"7400000400",x"3000000000",
		x"c000000232",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480040c0f",x"7400020400",x"3000000000",
		x"c000000233",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480020c0f",x"7400010400",x"3000000000",
		x"c000000234",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480060c0f",x"7400030400",x"3000000000",
		x"c000000235",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480010c0f",x"7400008400",x"3000000000",
		x"c000000236",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480050c0f",x"7400028400",x"3000000000",
		x"c000000237",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480030c0f",x"7400018400",x"3000000000",
		x"c000000238",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480070c0f",x"7400038400",x"3000000000",
		x"c000000239",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480008c0f",x"7400004400",x"3000000000",
		x"c00000023a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480048c0f",x"7400024400",x"3000000000",
		x"c00000023b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480028c0f",x"7400014400",x"3000000000",
		x"c00000023c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480068c0f",x"7400034400",x"3000000000",
		x"c00000023d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480018c0f",x"740000c400",x"3000000000",
		x"c00000023e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480058c0f",x"740002c400",x"3000000000",
		x"c00000023f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480038c0f",x"740001c400",x"3000000000",
		x"c000000240",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480078c0f",x"740003c400",x"3000000000",
		x"c000000241",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480004c0f",x"7400002400",x"3000000000",
		x"c000000242",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480044c0f",x"7400022400",x"3000000000",
		x"c000000243",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480024c0f",x"7400012400",x"3000000000",
		x"c000000244",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480064c0f",x"7400032400",x"3000000000",
		x"c000000245",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480014c0f",x"740000a400",x"3000000000",
		x"c000000246",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480054c0f",x"740002a400",x"3000000000",
		x"c000000247",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480034c0f",x"740001a400",x"3000000000",
		x"c000000248",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480074c0f",x"740003a400",x"3000000000",
		x"c000000249",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000cc0f",x"7400006400",x"3000000000",
		x"c00000024a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004cc0f",x"7400026400",x"3000000000",
		x"c00000024b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002cc0f",x"7400016400",x"3000000000",
		x"c00000024c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006cc0f",x"7400036400",x"3000000000",
		x"c00000024d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001cc0f",x"740000e400",x"3000000000",
		x"c00000024e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005cc0f",x"740002e400",x"3000000000",
		x"c00000024f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003cc0f",x"740001e400",x"3000000000",
		x"c000000250",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007cc0f",x"740003e400",x"3000000000",
		x"c000000251",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480002c0f",x"7400001400",x"3000000000",
		x"c000000252",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480042c0f",x"7400021400",x"3000000000",
		x"c000000253",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480022c0f",x"7400011400",x"3000000000",
		x"c000000254",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480062c0f",x"7400031400",x"3000000000",
		x"c000000255",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480012c0f",x"7400009400",x"3000000000",
		x"c000000256",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480052c0f",x"7400029400",x"3000000000",
		x"c000000257",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480032c0f",x"7400019400",x"3000000000",
		x"c000000258",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480072c0f",x"7400039400",x"3000000000",
		x"c000000259",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000ac0f",x"7400005400",x"3000000000",
		x"c00000025a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004ac0f",x"7400025400",x"3000000000",
		x"c00000025b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002ac0f",x"7400015400",x"3000000000",
		x"c00000025c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006ac0f",x"7400035400",x"3000000000",
		x"c00000025d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001ac0f",x"740000d400",x"3000000000",
		x"c00000025e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005ac0f",x"740002d400",x"3000000000",
		x"c00000025f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003ac0f",x"740001d400",x"3000000000",
		x"c000000260",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007ac0f",x"740003d400",x"3000000000",
		x"c000000261",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480006c0f",x"7400003400",x"3000000000",
		x"c000000262",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480046c0f",x"7400023400",x"3000000000",
		x"c000000263",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480026c0f",x"7400013400",x"3000000000",
		x"c000000264",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480066c0f",x"7400033400",x"3000000000",
		x"c000000265",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480016c0f",x"740000b400",x"3000000000",
		x"c000000266",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480056c0f",x"740002b400",x"3000000000",
		x"c000000267",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480036c0f",x"740001b400",x"3000000000",
		x"c000000268",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480076c0f",x"740003b400",x"3000000000",
		x"c000000269",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000ec0f",x"7400007400",x"3000000000",
		x"c00000026a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004ec0f",x"7400027400",x"3000000000",
		x"c00000026b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002ec0f",x"7400017400",x"3000000000",
		x"c00000026c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006ec0f",x"7400037400",x"3000000000",
		x"c00000026d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001ec0f",x"740000f400",x"3000000000",
		x"c00000026e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005ec0f",x"740002f400",x"3000000000",
		x"c00000026f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003ec0f",x"740001f400",x"3000000000",
		x"c000000270",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007ec0f",x"740003f400",x"3000000000",
		x"c000000271",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480001c0f",x"7400000c00",x"3000000000",
		x"c000000272",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480041c0f",x"7400020c00",x"3000000000",
		x"c000000273",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480021c0f",x"7400010c00",x"3000000000",
		x"c000000274",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480061c0f",x"7400030c00",x"3000000000",
		x"c000000275",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480011c0f",x"7400008c00",x"3000000000",
		x"c000000276",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480051c0f",x"7400028c00",x"3000000000",
		x"c000000277",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480031c0f",x"7400018c00",x"3000000000",
		x"c000000278",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480071c0f",x"7400038c00",x"3000000000",
		x"c000000279",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480009c0f",x"7400004c00",x"3000000000",
		x"c00000027a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480049c0f",x"7400024c00",x"3000000000",
		x"c00000027b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480029c0f",x"7400014c00",x"3000000000",
		x"c00000027c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480069c0f",x"7400034c00",x"3000000000",
		x"c00000027d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480019c0f",x"740000cc00",x"3000000000",
		x"c00000027e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480059c0f",x"740002cc00",x"3000000000",
		x"c00000027f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480039c0f",x"740001cc00",x"3000000000",
		x"c000000280",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480079c0f",x"740003cc00",x"3000000000",
		x"c000000281",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480005c0f",x"7400002c00",x"3000000000",
		x"c000000282",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480045c0f",x"7400022c00",x"3000000000",
		x"c000000283",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480025c0f",x"7400012c00",x"3000000000",
		x"c000000284",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480065c0f",x"7400032c00",x"3000000000",
		x"c000000285",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480015c0f",x"740000ac00",x"3000000000",
		x"c000000286",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480055c0f",x"740002ac00",x"3000000000",
		x"c000000287",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480035c0f",x"740001ac00",x"3000000000",
		x"c000000288",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480075c0f",x"740003ac00",x"3000000000",
		x"c000000289",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000dc0f",x"7400006c00",x"3000000000",
		x"c00000028a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004dc0f",x"7400026c00",x"3000000000",
		x"c00000028b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002dc0f",x"7400016c00",x"3000000000",
		x"c00000028c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006dc0f",x"7400036c00",x"3000000000",
		x"c00000028d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001dc0f",x"740000ec00",x"3000000000",
		x"c00000028e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005dc0f",x"740002ec00",x"3000000000",
		x"c00000028f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003dc0f",x"740001ec00",x"3000000000",
		x"c000000290",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007dc0f",x"740003ec00",x"3000000000",
		x"c000000291",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480003c0f",x"7400001c00",x"3000000000",
		x"c000000292",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480043c0f",x"7400021c00",x"3000000000",
		x"c000000293",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480023c0f",x"7400011c00",x"3000000000",
		x"c000000294",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480063c0f",x"7400031c00",x"3000000000",
		x"c000000295",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480013c0f",x"7400009c00",x"3000000000",
		x"c000000296",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480053c0f",x"7400029c00",x"3000000000",
		x"c000000297",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480033c0f",x"7400019c00",x"3000000000",
		x"c000000298",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480073c0f",x"7400039c00",x"3000000000",
		x"c000000299",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000bc0f",x"7400005c00",x"3000000000",
		x"c00000029a",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004bc0f",x"7400025c00",x"3000000000",
		x"c00000029b",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002bc0f",x"7400015c00",x"3000000000",
		x"c00000029c",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006bc0f",x"7400035c00",x"3000000000",
		x"c00000029d",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001bc0f",x"740000dc00",x"3000000000",
		x"c00000029e",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005bc0f",x"740002dc00",x"3000000000",
		x"c00000029f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003bc0f",x"740001dc00",x"3000000000",
		x"c0000002a0",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007bc0f",x"740003dc00",x"3000000000",
		x"c0000002a1",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480007c0f",x"7400003c00",x"3000000000",
		x"c0000002a2",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480047c0f",x"7400023c00",x"3000000000",
		x"c0000002a3",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480027c0f",x"7400013c00",x"3000000000",
		x"c0000002a4",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480067c0f",x"7400033c00",x"3000000000",
		x"c0000002a5",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480017c0f",x"740000bc00",x"3000000000",
		x"c0000002a6",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480057c0f",x"740002bc00",x"3000000000",
		x"c0000002a7",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480037c0f",x"740001bc00",x"3000000000",
		x"c0000002a8",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"4480077c0f",x"740003bc00",x"3000000000",
		x"c0000002a9",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448000fc0f",x"7400007c00",x"3000000000",
		x"c0000002aa",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448004fc0f",x"7400027c00",x"3000000000",
		x"c0000002ab",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448002fc0f",x"7400017c00",x"3000000000",
		x"c0000002ac",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448006fc0f",x"7400037c00",x"3000000000",
		x"c0000002ad",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448001fc0f",x"740000fc00",x"3000000000",
		x"c0000002ae",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448005fc0f",x"740002fc00",x"3000000000",
		x"c0000002af",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448003fc0f",x"740001fc00",x"3000000000",
		x"408000000f",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"3000000000",x"448007fc0f",x"740003fc00",x"3000000000"
	);
end ccsds_constants;

package body ccsds_constants is
	
end ccsds_constants;
