----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02.03.2021 10:35:20
-- Design Name: 
-- Module Name: constants - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package ccsds_test_constants is
	CONSTANT CONST_GOLDEN_NUM_S 	   	: integer := 0;
	CONSTANT CONST_GOLDEN_NUM_DRPSV 	: integer := 1;
	CONSTANT CONST_GOLDEN_NUM_PSV 		: integer := 2;
	CONSTANT CONST_GOLDEN_NUM_PR 		: integer := 3;
	CONSTANT CONST_GOLDEN_NUM_W			: integer := 4;
	CONSTANT CONST_GOLDEN_NUM_WUSE  	: integer := 5;
	CONSTANT CONST_GOLDEN_NUM_DRPE  	: integer := 6;
	CONSTANT CONST_GOLDEN_NUM_DRSR  	: integer := 7;
	CONSTANT CONST_GOLDEN_NUM_CQBC  	: integer := 8;
	CONSTANT CONST_GOLDEN_NUM_MEV 		: integer := 9;
	CONSTANT CONST_GOLDEN_NUM_HRPS   	: integer := 10;
	CONSTANT CONST_GOLDEN_NUM_PCD 		: integer := 11;
	CONSTANT CONST_GOLDEN_NUM_CLD 		: integer := 12;
	CONSTANT CONST_GOLDEN_NUM_NWD 		: integer := 13;
	CONSTANT CONST_GOLDEN_NUM_WD 		: integer := 14;
	CONSTANT CONST_GOLDEN_NUM_ND 		: integer := 15;
	CONSTANT CONST_GOLDEN_NUM_LS 		: integer := 16;
	CONSTANT CONST_GOLDEN_NUM_QI 		: integer := 17;
	CONSTANT CONST_GOLDEN_NUM_SR 		: integer := 18;
	CONSTANT CONST_GOLDEN_NUM_TS 		: integer := 19;
	CONSTANT CONST_GOLDEN_NUM_MQI 		: integer := 20;
	CONSTANT CONST_GOLDEN_NUM_ACC 		: integer := 21;
end ccsds_test_constants;

package body ccsds_test_constants is
	
end ccsds_test_constants;
