----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04.03.2021 12:38:18
-- Design Name: 
-- Module Name: ccsds_123b2_core - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.ccsds_constants.all;
use work.ccsds_data_structures.all;
use IEEE.NUMERIC_STD.ALL;
use work.am_data_types.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ccsds_123b2_core is
--	generic (
--		MAX_X_WIDTH: integer := 9;
--		MAX_Y_WIDTH: integer := 10;
--		MAX_Z_WIDTH: integer := 8;
--		MAX_T_WIDTH: integer := 19;
--		DATA_WIDTH: integer := CONST_MAX_D;
--		OUT_BYTES: integer := CONST_OUT_BYTES
--	);
--	port ( 

--	);
end ccsds_123b2_core;

architecture Behavioral of ccsds_123b2_core is
			
begin
	
end Behavioral;
