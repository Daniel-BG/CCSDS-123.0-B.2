----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02.03.2021 10:35:20
-- Design Name: 
-- Module Name: constants - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.ccsds_math_functions.all;

package ccsds_constants is
	--IMAGE CONSTANTS
	type local_sum_t is (WIDE_NEIGHBOR_ORIENTED, WIDE_COLUMN_ORIENTED);
	type relocation_mode_t is (VERTICAL_TO_DIAGONAL, DIAGONAL_TO_VERTICAL); 
	
	--OTHER CONSTANTS
	constant STDLV_ONE: std_logic_vector(0 downto 0) := "1";
	constant STDLV_ZERO: std_logic_vector(0 downto 0) := "0";
	
	--FIXED CONSTANTS
	constant CONST_TINC_MIN				: integer := 4;
	constant CONST_TINC_MAX				: integer := 11;
	constant CONST_TINC_BITS 			: integer := 4;
	constant CONST_VMIN					: integer := -6;
	constant CONST_VMAX					: integer := 9;
	constant CONST_VMINMAX_BITS 		: integer := 5;
	constant CONST_WEO_MIN				: integer := -6;
	constant CONST_WEO_MAX				: integer := 5;
	constant CONST_WEO_BITS 			: integer := 4;
	constant CONST_MAX_RES_VAL 			: integer := 4;
	constant CONST_DATA_WIDTH_MAX		: integer := 32;
	constant CONST_DATA_WIDTH_MIN		: integer := 2;
	constant CONST_OMEGA_WIDTH_MAX		: integer := 19;
	constant CONST_OMEGA_WIDTH_MIN		: integer := 4;
	constant CONST_WUSE_BITS 			: integer := 7;

	--CONSTANTS THAT CAN ALTER RESOURCE USE
	constant CONST_MAX_DATA_WIDTH		: integer := 16;				--maximum allowed bits for inputs (Can be set lower through cfg ports)
	constant CONST_MAX_OMEGA			: integer := 19;				--maximum allowed bits for weights (Can be set lower through cfg ports)
	constant CONST_MIN_OMEGA			: integer := 4;
	constant CONST_MAX_P				: integer := 3;					--maximum allowed bits for previous bands used in prediction
	constant CONST_MAX_BANDS			: integer := 256;				--maximum allowed size in the x direction (Can be set lower through cfg ports)
	constant CONST_MAX_LINES			: integer := 1024;				--maximum allowed size in the y direction (Can be set lower through cfg ports)
	constant CONST_MAX_SAMPLES			: integer := 512;  				--maximum allowed size in the z direction (Can be set lower through cfg ports)
	
	--DERIVED CONSTANTS
	constant CONST_MAX_SAMPLES_PER_BAND	: integer := CONST_MAX_SAMPLES * CONST_MAX_LINES;
	
	constant CONST_MAX_X_VALUE			: integer := CONST_MAX_SAMPLES - 1;	--maximum allowed size in the x direction (Can be set lower through cfg ports)
	constant CONST_MAX_Y_VALUE			: integer := CONST_MAX_LINES - 1;	--maximum allowed size in the y direction (Can be set lower through cfg ports)
	constant CONST_MAX_Z_VALUE			: integer := CONST_MAX_BANDS - 1;  	--maximum allowed size in the z direction (Can be set lower through cfg ports)
	constant CONST_MAX_T_VALUE			: integer := CONST_MAX_SAMPLES_PER_BAND - 1;
	
	constant CONST_ABS_ERR_BITS 		: integer := MIN(CONST_MAX_DATA_WIDTH - 1, 16); 
	constant CONST_REL_ERR_BITS 		: integer := MIN(CONST_MAX_DATA_WIDTH - 1, 16); 
	
	constant CONST_MAX_WEIGHT_BITS		: integer := CONST_MAX_OMEGA + 3;
	constant CONST_MAX_C				: integer := CONST_MAX_P + 3; --number of previous bands plus 3 (full pred mode)
	constant CONST_MAX_OMEGA_WIDTH_BITS	: integer := BITS(CONST_MAX_OMEGA);		
	constant CONST_MAX_DATA_WIDTH_BITS	: integer := BITS(CONST_MAX_DATA_WIDTH);	
	constant CONST_MAX_P_WIDTH_BITS  	: integer := BITS(CONST_MAX_P);
	constant CONST_MAX_C_BITS			: integer := BITS(CONST_MAX_C);
	
	constant CONST_MAX_X_VALUE_BITS		: integer := BITS(CONST_MAX_X_VALUE);
	constant CONST_MAX_Y_VALUE_BITS		: integer := BITS(CONST_MAX_Y_VALUE);
	constant CONST_MAX_Z_VALUE_BITS		: integer := BITS(CONST_MAX_Z_VALUE);
	constant CONST_MAX_T_VALUE_BITS		: integer := BITS(CONST_MAX_T_VALUE);
	
	constant CONST_MAX_BANDS_BITS		: integer := BITS(CONST_MAX_BANDS);
	constant CONST_MAX_LINES_BITS		: integer := BITS(CONST_MAX_LINES);
	constant CONST_MAX_SAMPLES_BITS		: integer := BITS(CONST_MAX_SAMPLES);
	
	constant CONST_CQBC_BITS			: integer := CONST_MAX_DATA_WIDTH;
	constant CONST_QI_BITS				: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_LSUM_BITS			: integer := CONST_MAX_DATA_WIDTH + 2;
	constant CONST_LDIF_BITS			: integer := CONST_MAX_DATA_WIDTH + 3;
	constant CONST_DRSR_BITS 			: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_DRPSV_BITS 			: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_DRPE_BITS 			: integer := CONST_MAX_DATA_WIDTH + 2;
	constant CONST_PR_BITS 				: integer := CONST_MAX_DATA_WIDTH + 1;
	
	constant CONST_MEV_BITS 			: integer := MAX(CONST_ABS_ERR_BITS, CONST_REL_ERR_BITS);
	constant CONST_PCLD_BITS 			: integer := CONST_MAX_WEIGHT_BITS + CONST_MAX_DATA_WIDTH + BITS(8*CONST_MAX_P + 19);
	constant CONST_HRPSV_BITS			: integer := CONST_MAX_OMEGA + 2 + CONST_MAX_DATA_WIDTH;
	
	constant CONST_RES_BITS				: integer := BITS(CONST_MAX_RES_VAL);
	constant CONST_DAMPING_BITS			: integer := CONST_MAX_RES_VAL;
	constant CONST_OFFSET_BITS			: integer := CONST_MAX_RES_VAL;
	
	constant CONST_DIFFVEC_BITS 		: integer := CONST_MAX_C * CONST_LDIF_BITS;
	constant CONST_CLDVEC_BITS 			: integer := CONST_MAX_P * CONST_LDIF_BITS;
	constant CONST_DIRDIFFVEC_BITS		: integer := 3 * CONST_LDIF_BITS;
	constant CONST_WEIGHTVEC_BITS		: integer := CONST_MAX_C * CONST_MAX_WEIGHT_BITS;
	
	constant CONST_W_UPDATE_BITS		: integer := CONST_LDIF_BITS - CONST_VMIN - CONST_WEO_MIN - CONST_DATA_WIDTH_MIN + CONST_OMEGA_WIDTH_MAX; --should be 64
	
	constant CONST_THETA_BITS			: integer := CONST_MAX_DATA_WIDTH;
	constant CONST_MQI_BITS				: integer := CONST_MAX_DATA_WIDTH;
	
	--ENCODER OUTPUT CONSTANTS
	constant CONST_OUTPUT_CODE_LENGTH 	: integer := 64;
	constant CONST_OUTPUT_CODE_LENGTH_BITS: integer := 7;
	
	--ENCODER CONSTANTS
	constant CONST_MIN_GAMMA_ZERO		: integer := 1;
	constant CONST_MAX_GAMMA_ZERO		: integer := 8;
	constant CONST_MAX_GAMMA_STAR		: integer := 11;
	constant CONST_MAX_GAMMA_STAR_BITS	: integer := BITS(CONST_MAX_GAMMA_STAR);
	constant CONST_MAX_COUNTER_BITS 	: integer := CONST_MAX_GAMMA_STAR;
	constant CONST_MAX_ACC_BITS			: integer := CONST_MAX_GAMMA_STAR + CONST_MAX_DATA_WIDTH;
	constant CONST_MAX_HR_ACC_BITS		: integer := CONST_MAX_ACC_BITS + 2;
	constant CONST_MAX_K				: integer := CONST_MAX_DATA_WIDTH - 2;
	constant CONST_MAX_K_BITS			: integer := BITS(CONST_MAX_K);
	constant CONST_U_MAX_MIN			: integer := 8;
	constant CONST_U_MAX_MAX			: integer := 32;
	constant CONST_U_MAX_BITS			: integer := BITS(CONST_U_MAX_MAX);
	
	constant CONST_MAX_CODE_LENGTH		: integer := CONST_U_MAX_MAX + CONST_MAX_DATA_WIDTH;
	constant CONST_MAX_CODE_LENGTH_BITS : integer := BITS(CONST_MAX_CODE_LENGTH);
	
	--HYBRID ENCODER SPECIFIC CONSTANTS
	constant CONST_LE_TABLE_COUNT: integer := 16;
	constant CONST_CODE_INDEX_BITS: integer := bits(CONST_LE_TABLE_COUNT - 1);
	
	constant CONST_MAX_THRESHOLD_VALUE_BITS : integer := 19;
	subtype threshold_value_t is std_logic_vector (CONST_MAX_THRESHOLD_VALUE_BITS - 1 downto 0);
    type threshold_table_t is array (0 to CONST_LE_TABLE_COUNT - 1) of threshold_value_t;

    constant CONST_THRESHOLD_TABLE : threshold_table_t := (
		"100" & x"A0E8",
		"011" & x"707C",
		"010" & x"8C43",
		"001" & x"F6A0",
		"001" & x"756D",
		"001" & x"1026",
		"000" & x"C5F6",
		"000" & x"8852",
		"000" & x"5B23",
		"000" & x"3A57",
		"000" & x"2442",
		"000" & x"1586",
		"000" & x"0C7B",
		"000" & x"0788",
		"000" & x"0458",
		"000" & x"0198"
	);
	
	constant CONST_INPUT_SYMBOL_AMOUNT: integer := 15;
	constant CONST_INPUT_SYMBOL_BITS: integer := bits(CONST_INPUT_SYMBOL_AMOUNT - 1);
	constant CONST_INPUT_SYMBOL_X	 : std_logic_vector := std_logic_vector(to_unsigned(13, CONST_INPUT_SYMBOL_BITS)); --"1101";
	constant CONST_INPUT_SYMBOL_FLUSH: std_logic_vector := std_logic_vector(to_unsigned(14, CONST_INPUT_SYMBOL_BITS)); --"1110";
	
	type input_symbol_limit_t is array (0 to CONST_LE_TABLE_COUNT - 1) of std_logic_vector(CONST_INPUT_SYMBOL_BITS - 1 downto 0);
	constant CONST_INPUT_SYMBOL_LIMIT : input_symbol_limit_t := (
		x"C", x"A", x"8", x"6",
		x"6", x"4", x"4", x"4",
		x"2", x"2", x"2", x"2",
		x"2", x"2", x"2", x"0"		
	);
	
	constant CONST_CODEWORD_BITS: integer := 21;
	constant CONST_CODEWORD_LENGTH_BITS: integer := 5;
	
	constant CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT: integer := 688;
	constant CONST_LOW_ENTROPY_CODING_TABLE_ADDRESS_BITS: integer := bits(CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT);
	
	constant CONST_LOW_ENTROPY_TABLE_ENTRY_BITS: integer := 32;

	type table_rom_t_v2 is array(0 to CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT*16 - 1) of std_logic_vector(CONST_LOW_ENTROPY_TABLE_ENTRY_BITS - 1 downto 0);
	constant CONST_LOW_ENTROPY_CODING_TABLE_V2: table_rom_t_v2 := (
		x"40000010",x"c0600000",x"c0600004",x"c0600002",x"40000011",x"c0800006",x"c080000e",x"40000012",x"40000013",x"c0a00001",x"c0a00011",x"c0c00005",x"c0c00025",x"c0a00009",x"f0200000",x"b0000000",
		x"40000014",x"40000015",x"40000016",x"c0600000",x"c0600004",x"c0800002",x"c080000a",x"c0a00006",x"c0a00016",x"c0c0000d",x"40000017",x"b0000000",x"b0000000",x"c0c0002d",x"f0200000",x"b0000000",
		x"c0400000",x"40000018",x"40000019",x"c0600002",x"c0600006",x"4000001a",x"4000001b",x"c0c00019",x"c0c00039",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c0c00005",x"f0200000",x"b0000000",
		x"4000001c",x"c0400000",x"4000001d",x"4000001e",x"4000001f",x"c0a0000e",x"40000020",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c0c00005",x"f0200000",x"b0000000",
		x"40000021",x"c0400000",x"c0400002",x"c0800001",x"c0800009",x"c0e00013",x"c0e00053",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1000027",x"f0200000",x"b0000000",
		x"c0200000",x"c0400001",x"40000022",x"c0a00003",x"c0a00013",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c0e0001b",x"f0200000",x"b0000000",
		x"40000023",x"40000024",x"40000025",x"40000026",x"c0e0000b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120006f",x"f0400000",x"b0000000",
		x"40000027",x"40000028",x"c0600001",x"40000029",x"c12000ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c14001bf",x"f0200000",x"b0000000",
		x"4000002a",x"4000002b",x"4000002c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120006f",x"f0400000",x"b0000000",
		x"4000002d",x"c0800002",x"c080000a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c140005f",x"f0600000",x"b0000000",
		x"4000002e",x"4000002f",x"c0a00001",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18005ff",x"f0600000",x"b0000000",
		x"40000030",x"c0a00001",x"40000031",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c00bff",x"f0800000",x"b0000000",
		x"40000032",x"c0c00001",x"c0c00021",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e01bff",x"f0800000",x"b0000000",
		x"40000033",x"40000034",x"c0e00001",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e003ff",x"f0a00000",x"b0000000",
		x"40000035",x"c1000001",x"c1000081",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20003ff",x"f0c00000",x"b0000000",
		x"40000036",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200001",x"f1000000",x"b0000000",
		x"c0a00019",x"40000037",x"40000038",x"c0c00015",x"c0c00035",x"c0c0000d",x"c0c0002d",x"c0e00013",x"c0e00053",x"c100003b",x"c10000bb",x"c120000f",x"c120010f",x"c100007b",x"f0400001",x"b0000000",
		x"c0c0001d",x"c0c0003d",x"c0c00003",x"c0c00023",x"40000039",x"c0e00033",x"c0e00073",x"c10000fb",x"c1000007",x"c120008f",x"c120018f",x"c120004f",x"c120014f",x"c1000087",x"f0600003",x"b0000000",
		x"c0e0000b",x"c0e0004b",x"c0e0002b",x"c1000047",x"c10000c7",x"c1000027",x"c10000a7",x"c12000cf",x"c12001cf",x"c140015f",x"c140035f",x"c160007f",x"c160047f",x"c14000df",x"f0a00007",x"b0000000",
		x"c0e0006b",x"c0e0001b",x"c0e0005b",x"c1000067",x"c10000e7",x"c1000017",x"c1000097",x"c120002f",x"c120012f",x"c14002df",x"c14001df",x"c160027f",x"c160067f",x"c14003df",x"f0a00017",x"b0000000",
		x"4000003a",x"c0a0000e",x"c0a0001e",x"4000003b",x"4000003c",x"c0c0001d",x"c0c0003d",x"c0e00013",x"c0e00053",x"c12000e7",x"c12001e7",x"b0000000",x"b0000000",x"c100002b",x"f0600001",x"b0000000",
		x"c0a00001",x"c0a00011",x"c0a00009",x"4000003d",x"c0c00003",x"4000003e",x"4000003f",x"c10000ab",x"c100006b",x"c1200017",x"c1200117",x"b0000000",x"b0000000",x"c1200097",x"f0600005",x"b0000000",
		x"c0a00019",x"c0a00005",x"c0a00015",x"40000040",x"c0c00023",x"40000041",x"c0e00033",x"c10000eb",x"c100001b",x"c1200197",x"c1200057",x"b0000000",x"b0000000",x"c1200157",x"f0600003",x"b0000000",
		x"c12000d7",x"c12001d7",x"c1200037",x"c14001ef",x"c14003ef",x"c140001f",x"c140021f",x"c160023f",x"c180017f",x"c1a00dff",x"c1a01dff",x"b0000000",x"b0000000",x"c180097f",x"f0e0001f",x"b0000000",
		x"c0800001",x"40000042",x"40000043",x"40000044",x"40000045",x"c0e00035",x"c0e00075",x"c100006b",x"c12000f7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001f7",x"f0600001",x"b0000000",
		x"40000046",x"40000047",x"c0a00009",x"40000048",x"40000049",x"c0e0000d",x"c0e0004d",x"c10000eb",x"c120000f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120010f",x"f0600005",x"b0000000",
		x"c0c00025",x"c0e0002d",x"c0e0006d",x"c100001b",x"c100009b",x"c120008f",x"c120018f",x"c16000bf",x"c16004bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16002bf",x"f0a00003",x"b0000000",
		x"c0e0001d",x"c0e0005d",x"c0e0003d",x"c100005b",x"c10000db",x"c120004f",x"c120014f",x"c16006bf",x"c16001bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16005bf",x"f0a00013",x"b0000000",
		x"4000004a",x"c0800002",x"c080000a",x"c0a0001e",x"c0a00001",x"c0e0002d",x"c0e0006d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c100006b",x"f0600001",x"b0000000",
		x"c0800006",x"4000004b",x"4000004c",x"4000004d",x"c0c00025",x"c10000eb",x"c100001b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c100009b",x"f0600005",x"b0000000",
		x"c0a00011",x"4000004e",x"4000004f",x"c0e0001d",x"c0e0005d",x"c1200077",x"c1200177",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000f7",x"f0800003",x"b0000000",
		x"c0a00009",x"40000050",x"c0c00015",x"c0e0003d",x"c0e0007d",x"c12001f7",x"c120000f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c14000df",x"f0a00007",x"b0000000",
		x"c0e00003",x"c100005b",x"c10000db",x"c120010f",x"c120008f",x"c16002bf",x"c16006bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18002ff",x"f0e0000f",x"b0000000",
		x"40000051",x"40000052",x"40000053",x"40000054",x"40000055",x"c10000a7",x"c1000067",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000ef",x"f0400001",x"b0000000",
		x"40000056",x"40000057",x"40000058",x"c0e0005b",x"40000059",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000b7",x"f0600001",x"b0000000",
		x"4000005a",x"c0600000",x"4000005b",x"c0e0004b",x"c0e0002b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120016f",x"f0400002",x"b0000000",
		x"c0600004",x"4000005c",x"c0a00009",x"c12000ef",x"c12001ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16001bf",x"f0800005",x"b0000000",
		x"4000005d",x"c0a00019",x"c0a00005",x"c120001f",x"c120011f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16005bf",x"f080000d",x"b0000000",
		x"c0e0006b",x"c120009f",x"c120019f",x"c1a005ff",x"c1a015ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e03fff",x"f100007f",x"b0000000",
		x"c0200000",x"4000005e",x"4000005f",x"c12001ef",x"c120001f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160027f",x"f0400001",x"b0000000",
		x"40000060",x"40000061",x"c0c0000b",x"c160067f",x"c160017f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a003ff",x"f0800003",x"b0000000",
		x"c120011f",x"c160057f",x"c160037f",x"c2001fff",x"c220bfff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c241ffff",x"f12000ff",x"b0000000",
		x"40000062",x"40000063",x"c0800004",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120016f",x"f0600002",x"b0000000",
		x"40000064",x"40000065",x"c0e0001b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18001ff",x"f0c00007",x"b0000000",
		x"40000066",x"40000067",x"c0e0005b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18009ff",x"f0c00027",x"b0000000",
		x"40000068",x"c0800006",x"40000069",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16000ff",x"f0600004",x"b0000000",
		x"4000006a",x"4000006b",x"c0a00011",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800dff",x"f0600004",x"b0000000",
		x"4000006c",x"c120002f",x"c14001af",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2201fff",x"f100000f",x"b0000000",
		x"4000006d",x"4000006e",x"4000006f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c02bff",x"f0800008",x"b0000000",
		x"40000070",x"c160005f",x"c160045f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2837fff",x"f14000df",x"b0000000",
		x"40000071",x"c0c00011",x"40000072",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e05bff",x"f0800008",x"b0000000",
		x"40000073",x"c0e00041",x"c0e00021",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e043ff",x"f0a00010",x"b0000000",
		x"40000074",x"c18001ff",x"c18009ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c241ffff",x"f100007f",x"b0000000",
		x"40000075",x"c1000041",x"c10000c1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20083ff",x"f0c00020",x"b0000000",
		x"40000076",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200101",x"f1000080",x"b0000000",
		x"c1000057",x"c10000d7",x"c1000037",x"c12000af",x"c12001af",x"c120006f",x"c120016f",x"c140003f",x"c140023f",x"c160017f",x"c160057f",x"c18001ff",x"c18009ff",x"c160037f",x"f0a0000f",x"b0000000",
		x"c10000b7",x"c1000077",x"c10000f7",x"c12000ef",x"c12001ef",x"c120001f",x"c120011f",x"c140013f",x"c140033f",x"c160077f",x"c16000ff",x"c18005ff",x"c1800dff",x"c16004ff",x"f0c0001f",x"b0000000",
		x"c120009f",x"c120019f",x"c120005f",x"c14000bf",x"c14002bf",x"c14001bf",x"c14003bf",x"c16002ff",x"c16006ff",x"c18003ff",x"c1800bff",x"c1a00fff",x"c1a01fff",x"c18007ff",x"f0c0003f",x"b0000000",
		x"c0e00073",x"c0e0000b",x"c0e0004b",x"c100009b",x"c100005b",x"c1200137",x"c12000b7",x"c140011f",x"c140031f",x"c160063f",x"c160013f",x"b0000000",x"b0000000",x"c160053f",x"f0a00007",x"b0000000",
		x"c10000db",x"c100003b",x"c10000bb",x"c12001b7",x"c1200077",x"c1200177",x"c12000f7",x"c140009f",x"c160033f",x"c180057f",x"c1800d7f",x"b0000000",x"b0000000",x"c160073f",x"f0c00017",x"b0000000",
		x"c100007b",x"c10000fb",x"c1000007",x"c12001f7",x"c120000f",x"c120010f",x"c140029f",x"c16000bf",x"c16004bf",x"c180037f",x"c1800b7f",x"b0000000",x"b0000000",x"c16002bf",x"f0c00037",x"b0000000",
		x"c1000087",x"c1000047",x"c10000c7",x"c120008f",x"c120018f",x"c140019f",x"c140039f",x"c16006bf",x"c16001bf",x"c180077f",x"c1800f7f",x"b0000000",x"b0000000",x"c18000ff",x"f0c0000f",x"b0000000",
		x"c120004f",x"c120014f",x"c12000cf",x"c140005f",x"c140025f",x"c140015f",x"c16005bf",x"c18008ff",x"c18004ff",x"c1a003ff",x"c1a013ff",x"b0000000",x"b0000000",x"c1800cff",x"f0e0005f",x"b0000000",
		x"c12001cf",x"c120002f",x"c120012f",x"c140035f",x"c14000df",x"c16003bf",x"c16007bf",x"c18002ff",x"c1800aff",x"c1a00bff",x"c1a01bff",x"b0000000",x"b0000000",x"c1a007ff",x"f0e0003f",x"b0000000",
		x"c1000027",x"c10000a7",x"c1000067",x"c12000af",x"c12001af",x"c14002df",x"c14001df",x"c160007f",x"c160047f",x"c18006ff",x"c1800eff",x"b0000000",x"b0000000",x"c18001ff",x"f0c0002f",x"b0000000",
		x"c120006f",x"c120016f",x"c12000ef",x"c14003df",x"c140003f",x"c160027f",x"c160067f",x"c18009ff",x"c18005ff",x"c1a017ff",x"c1a00fff",x"b0000000",x"b0000000",x"c1a01fff",x"f0e0007f",x"b0000000",
		x"c0e0007d",x"c0e00003",x"c0e00043",x"c100003b",x"c10000bb",x"c12000cf",x"c12001cf",x"c16003bf",x"c16007bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160007f",x"f0a0000b",x"b0000000",
		x"c0e00023",x"c0e00063",x"c0e00013",x"c100007b",x"c10000fb",x"c120002f",x"c120012f",x"c160047f",x"c160027f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160067f",x"f0a0001b",x"b0000000",
		x"c0e00053",x"c1000007",x"c1000087",x"c12000af",x"c12001af",x"c14000df",x"c14002df",x"c18002ff",x"c1800aff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18006ff",x"f0c0000f",x"b0000000",
		x"c1000047",x"c10000c7",x"c1000027",x"c120006f",x"c120016f",x"c14001df",x"c14003df",x"c1800eff",x"c18001ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18009ff",x"f0c0002f",x"b0000000",
		x"c0c00015",x"c0e00033",x"c0e00073",x"c10000a7",x"c1000067",x"c12000ef",x"c12001ef",x"c160017f",x"c160057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160037f",x"f0a00007",x"b0000000",
		x"c0e0000b",x"c0e0004b",x"c0e0002b",x"c10000e7",x"c1000017",x"c120001f",x"c120011f",x"c160077f",x"c16000ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16004ff",x"f0a00017",x"b0000000",
		x"c1000097",x"c1000057",x"c10000d7",x"c120009f",x"c120019f",x"c140003f",x"c140023f",x"c18005ff",x"c1800dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18003ff",x"f0c0001f",x"b0000000",
		x"c1000037",x"c10000b7",x"c1000077",x"c120005f",x"c120015f",x"c140013f",x"c140033f",x"c1800bff",x"c18007ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800fff",x"f0c0003f",x"b0000000",
		x"c0a00019",x"40000077",x"40000078",x"c0e00043",x"c0e00023",x"c120018f",x"c120004f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120014f",x"f080000b",x"b0000000",
		x"c0c00035",x"40000079",x"c0e00063",x"c100003b",x"c10000bb",x"c14002df",x"c14001df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16001bf",x"f0c00017",x"b0000000",
		x"c0c0000d",x"4000007a",x"c0e00013",x"c100007b",x"c10000fb",x"c14003df",x"c140003f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16005bf",x"f0c00037",x"b0000000",
		x"c0e00053",x"c1000007",x"c1000087",x"c12000cf",x"c12001cf",x"c16003bf",x"c16007bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800aff",x"f0e0004f",x"b0000000",
		x"c0e00033",x"c1000047",x"c10000c7",x"c120002f",x"c120012f",x"c160007f",x"c160047f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18006ff",x"f0e0002f",x"b0000000",
		x"c0e00073",x"c1000027",x"c10000a7",x"c12000af",x"c12001af",x"c160027f",x"c160067f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800eff",x"f0e0006f",x"b0000000",
		x"c0e0000b",x"c1000067",x"c10000e7",x"c120006f",x"c120016f",x"c160017f",x"c160057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18001ff",x"f0e0001f",x"b0000000",
		x"c0800005",x"4000007b",x"c0a0000d",x"c0e00033",x"c0e00073",x"c12001ef",x"c140015f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c140035f",x"f0800003",x"b0000000",
		x"4000007c",x"4000007d",x"4000007e",x"c10000e7",x"c1000017",x"c14000df",x"c14002df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160017f",x"f080000b",x"b0000000",
		x"c0a0001d",x"4000007f",x"40000080",x"c1000097",x"c1000057",x"c14001df",x"c160057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160037f",x"f0a00007",x"b0000000",
		x"c0e0000b",x"c10000d7",x"c1000037",x"c120001f",x"c14003df",x"c180077f",x"c1800f7f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a005ff",x"f0c00017",x"b0000000",
		x"c0e0004b",x"c10000b7",x"c1000077",x"c140003f",x"c140023f",x"c18000ff",x"c1a015ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00dff",x"f0e0001f",x"b0000000",
		x"40000081",x"40000082",x"40000083",x"c100007b",x"c12001b7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c140019f",x"f0600005",x"b0000000",
		x"40000084",x"40000085",x"40000086",x"c140039f",x"c140005f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16000bf",x"f0a00003",x"b0000000",
		x"40000087",x"40000088",x"c0e0003b",x"c140025f",x"c140015f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c180027f",x"f0a00013",x"b0000000",
		x"c1200077",x"c140035f",x"c14000df",x"c1a00eff",x"c1a01eff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c00bff",x"f100003f",x"b0000000",
		x"40000089",x"4000008a",x"c0800006",x"c1000057",x"c10000d7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c140003f",x"f0600001",x"b0000000",
		x"c080000e",x"4000008b",x"c0c0000d",x"c140023f",x"c140013f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c180037f",x"f0a0000b",x"b0000000",
		x"4000008c",x"c0e0001b",x"c0e0005b",x"c16003bf",x"c1800b7f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00dff",x"f0c00007",x"b0000000",
		x"c0800001",x"4000008d",x"c0c0002d",x"c140033f",x"c14000bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c180077f",x"f0a0001b",x"b0000000",
		x"4000008e",x"c0c0002b",x"c0c0001b",x"c18004ff",x"c1800cff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c013ff",x"f0a0000b",x"b0000000",
		x"c0800005",x"c0c0003b",x"4000008f",x"c18002ff",x"c1800aff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c033ff",x"f0a0001b",x"b0000000",
		x"40000090",x"c0c00007",x"c0c00027",x"c18006ff",x"c1800eff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c00bff",x"f0a00007",x"b0000000",
		x"c0c00017",x"c100006f",x"40000091",x"c1c02bff",x"c1c01bff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2009fff",x"f0e0001f",x"b0000000",
		x"40000092",x"c080000c",x"c0800002",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c140003f",x"f0600006",x"b0000000",
		x"c080000a",x"c0e0003b",x"c0e0007b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a003ff",x"f0c00017",x"b0000000",
		x"c0800006",x"c0e00007",x"c0e00047",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18005ff",x"f0c00037",x"b0000000",
		x"c0e00027",x"c140023f",x"c140013f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e02fff",x"f120007f",x"b0000000",
		x"c080000e",x"c0e00067",x"c0e00017",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a013ff",x"f0e0000f",x"b0000000",
		x"c0e00057",x"c140033f",x"c14000bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2007fff",x"f14001ff",x"b0000000",
		x"40000093",x"40000094",x"40000095",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16004ff",x"f0600002",x"b0000000",
		x"40000096",x"c1000017",x"c12000f7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e007ff",x"f0e00007",x"b0000000",
		x"40000097",x"40000098",x"c0a00009",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a003ff",x"f0600002",x"b0000000",
		x"40000099",x"c120012f",x"c14003af",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2211fff",x"f100008f",x"b0000000",
		x"4000009a",x"c12000af",x"c140006f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2209fff",x"f100004f",x"b0000000",
		x"4000009b",x"4000009c",x"c0c00011",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c01bff",x"f0800004",x"b0000000",
		x"4000009d",x"c160025f",x"c160065f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2607fff",x"f120001f",x"b0000000",
		x"c0c00031",x"c160015f",x"c160055f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28b7fff",x"f14002df",x"b0000000",
		x"c0c00009",x"c160035f",x"c160075f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2877fff",x"f14001df",x"b0000000",
		x"4000009e",x"c0c00031",x"4000009f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e03bff",x"f0800004",x"b0000000",
		x"400000a0",x"c18000ff",x"c1a009ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c281ffff",x"f120003f",x"b0000000",
		x"400000a1",x"c0e00061",x"c0e00011",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e023ff",x"f0a00008",x"b0000000",
		x"c0e00051",x"c18005ff",x"c1800dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c243ffff",x"f10000ff",x"b0000000",
		x"400000a2",x"c1000021",x"c10000a1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20043ff",x"f0c00010",x"b0000000",
		x"400000a3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200081",x"f1000040",x"b0000000",
		x"c0e0004b",x"c1000017",x"c1000097",x"c12000ef",x"c12001ef",x"c160037f",x"c160077f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18009ff",x"f0e0005f",x"b0000000",
		x"c0e0002b",x"c1000057",x"c10000d7",x"c120001f",x"c120011f",x"c16000ff",x"c16004ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18005ff",x"f0e0003f",x"b0000000",
		x"c1000037",x"c120009f",x"c120019f",x"c140023f",x"c140013f",x"c1800dff",x"c18003ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00fff",x"f100007f",x"b0000000",
		x"c10000b7",x"c120005f",x"c120015f",x"c140033f",x"c14000bf",x"c1800bff",x"c18007ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a01fff",x"f10000ff",x"b0000000",
		x"c0c00003",x"c0e0002b",x"c0e0006b",x"c120011f",x"c120009f",x"c18008ff",x"c18004ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800cff",x"f0c00037",x"b0000000",
		x"c0c00023",x"c0e0001b",x"c0e0005b",x"c120019f",x"c120005f",x"c18002ff",x"c1800aff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18006ff",x"f0c0000f",x"b0000000",
		x"c0e0003b",x"c10000f7",x"c100000f",x"c140013f",x"c140033f",x"c1800eff",x"c1a01dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a003ff",x"f0c0002f",x"b0000000",
		x"c0e0007b",x"c100008f",x"c100004f",x"c14000bf",x"c14002bf",x"c18001ff",x"c1a013ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00bff",x"f0e0005f",x"b0000000",
		x"c0e00007",x"c10000cf",x"c100002f",x"c14001bf",x"c14003bf",x"c18009ff",x"c1a01bff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a007ff",x"f0e0003f",x"b0000000",
		x"c0e00047",x"c10000af",x"c100006f",x"c140007f",x"c140027f",x"c1a017ff",x"c1a00fff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a01fff",x"f0e0007f",x"b0000000",
		x"c0a0000b",x"400000a4",x"400000a5",x"c1200177",x"c14002df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16004bf",x"f0a0000b",x"b0000000",
		x"400000a6",x"c10000fb",x"c1000007",x"c16002bf",x"c16006bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a001ff",x"f0c0001b",x"b0000000",
		x"400000a7",x"c1000087",x"c1000047",x"c16001bf",x"c16005bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a011ff",x"f0c0003b",x"b0000000",
		x"400000a8",x"c10000c7",x"c1000027",x"c16003bf",x"c16007bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a009ff",x"f0c00007",x"b0000000",
		x"c10000a7",x"c12000f7",x"c12001f7",x"c1800a7f",x"c180067f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c02bff",x"f0e00037",x"b0000000",
		x"c1000067",x"c120000f",x"c120010f",x"c1800e7f",x"c180017f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c01bff",x"f0e00077",x"b0000000",
		x"400000a9",x"c10000e7",x"c1000017",x"c160007f",x"c160047f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a019ff",x"f0c00027",x"b0000000",
		x"c1000097",x"c120008f",x"c120018f",x"c180097f",x"c180057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c03bff",x"f0e0000f",x"b0000000",
		x"c0600002",x"400000aa",x"400000ab",x"c120005f",x"c120015f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16007bf",x"f0800003",x"b0000000",
		x"400000ac",x"c0c0001d",x"c0c0003d",x"c14002bf",x"c160007f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a01dff",x"f0c00027",x"b0000000",
		x"c0c00003",x"c1000037",x"c10000b7",x"c1800f7f",x"c18000ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c017ff",x"f0e0002f",x"b0000000",
		x"c0c00023",x"c1000077",x"c10000f7",x"c18008ff",x"c18004ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c037ff",x"f0e0006f",x"b0000000",
		x"400000ad",x"c100000f",x"c100008f",x"c1800cff",x"c18002ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c00fff",x"f0e0001f",x"b0000000",
		x"c080000d",x"400000ae",x"400000af",x"c18001ff",x"c18009ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c03bff",x"f0a00017",x"b0000000",
		x"c0e00037",x"c120009f",x"c120019f",x"c1e027ff",x"c1e067ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2005fff",x"f100005f",x"b0000000",
		x"c0800003",x"400000b0",x"400000b1",x"c18005ff",x"c1800dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c007ff",x"f0a0000f",x"b0000000",
		x"c120005f",x"c160077f",x"c16000ff",x"c200dfff",x"c221bfff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c243ffff",x"f12001ff",x"b0000000",
		x"400000b2",x"c0800001",x"400000b3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c14002bf",x"f0600001",x"b0000000",
		x"400000b4",x"400000b5",x"400000b6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16002ff",x"f0600006",x"b0000000",
		x"400000b7",x"c1000097",x"c1000057",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e047ff",x"f0e00047",x"b0000000",
		x"400000b8",x"c10000d7",x"c12001f7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e027ff",x"f0e00027",x"b0000000",
		x"400000b9",x"c1000037",x"c120000f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e067ff",x"f0e00067",x"b0000000",
		x"400000ba",x"c0a00019",x"c0a00005",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a013ff",x"f0600006",x"b0000000",
		x"c0a00015",x"c140026f",x"c140016f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2219fff",x"f10000cf",x"b0000000",
		x"c0a0000d",x"c140036f",x"c14000ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2205fff",x"f100002f",x"b0000000",
		x"c0a0001d",x"c14002ef",x"c14001ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2215fff",x"f10000af",x"b0000000",
		x"400000bb",x"400000bc",x"c0c00029",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c03bff",x"f080000c",x"b0000000",
		x"400000bd",x"c16000df",x"c16004df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2647fff",x"f120011f",x"b0000000",
		x"400000be",x"c16002df",x"c16006df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2627fff",x"f120009f",x"b0000000",
		x"400000bf",x"c0c00009",x"400000c0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e07bff",x"f080000c",x"b0000000",
		x"400000c1",x"c18008ff",x"c1a019ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c289ffff",x"f120013f",x"b0000000",
		x"400000c2",x"c18004ff",x"c1a005ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c285ffff",x"f12000bf",x"b0000000",
		x"400000c3",x"c0e00031",x"c0e00071",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e063ff",x"f0a00018",x"b0000000",
		x"400000c4",x"c1000061",x"c10000e1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200c3ff",x"f0c00030",x"b0000000",
		x"400000c5",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200181",x"f10000c0",x"b0000000",
		x"400000c6",x"c120004f",x"c120014f",x"c1800d7f",x"c180037f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c007ff",x"f0e0004f",x"b0000000",
		x"c1000057",x"c12000cf",x"c12001cf",x"c1800b7f",x"c180077f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c027ff",x"f0e0002f",x"b0000000",
		x"400000c7",x"c120002f",x"c120012f",x"c1800f7f",x"c18000ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c017ff",x"f0e0006f",x"b0000000",
		x"c10000d7",x"c12000af",x"c12001af",x"c18008ff",x"c18004ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c037ff",x"f0e0001f",x"b0000000",
		x"400000c8",x"c120006f",x"c120016f",x"c1800cff",x"c18002ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c00fff",x"f0c00017",x"b0000000",
		x"c1000037",x"c12000ef",x"c12001ef",x"c1800aff",x"c18006ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c02fff",x"f0e0005f",x"b0000000",
		x"400000c9",x"c0e0003b",x"c0e0007b",x"c160047f",x"c160027f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a003ff",x"f0c00017",x"b0000000",
		x"400000ca",x"c0e00007",x"c0e00047",x"c160067f",x"c1800aff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a013ff",x"f0c00037",x"b0000000",
		x"c0a00015",x"c0e00027",x"c0e00067",x"c160017f",x"c160057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00bff",x"f0c0000f",x"b0000000",
		x"c0e00017",x"c12000df",x"c12001df",x"c1a01bff",x"c1a007ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e07fff",x"f10000ff",x"b0000000",
		x"c0e00077",x"c120015f",x"c12000df",x"c1e017ff",x"c1e057ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2207fff",x"f10000df",x"b0000000",
		x"c0e0000f",x"c12001df",x"c14003bf",x"c1e037ff",x"c1e077ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2217fff",x"f100003f",x"b0000000",
		x"c0e0004f",x"c120003f",x"c120013f",x"c1e00fff",x"c1e04fff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2003fff",x"f10000bf",x"b0000000",
		x"c0e0002f",x"c12000bf",x"c140007f",x"c1e02fff",x"c1e06fff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220ffff",x"f100007f",x"b0000000",
		x"400000cb",x"400000cc",x"400000cd",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c14001bf",x"f0800005",x"b0000000",
		x"400000ce",x"400000cf",x"c1000077",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00bff",x"f0e0004f",x"b0000000",
		x"400000d0",x"400000d1",x"c0a0000e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16006ff",x"f0800001",x"b0000000",
		x"400000d2",x"c10000b7",x"c120010f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e017ff",x"f0e00017",x"b0000000",
		x"c0a0001e",x"c120008f",x"c120018f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2002fff",x"f100004f",x"b0000000",
		x"400000d3",x"c1000077",x"c120004f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e057ff",x"f0e00057",x"b0000000",
		x"c0a00001",x"c120014f",x"c12000cf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200afff",x"f10000cf",x"b0000000",
		x"c0a00011",x"c12001cf",x"c120002f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e037ff",x"f100002f",x"b0000000",
		x"400000d4",x"c0a00003",x"400000d5",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00bff",x"f0600001",x"b0000000",
		x"400000d6",x"400000d7",x"c0c00019",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c007ff",x"f0800002",x"b0000000",
		x"400000d8",x"c16001df",x"c16005df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2667fff",x"f120019f",x"b0000000",
		x"400000d9",x"c16003df",x"c16007df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2617fff",x"f120005f",x"b0000000",
		x"400000da",x"c160003f",x"c160043f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2657fff",x"f120015f",x"b0000000",
		x"400000db",x"c0c00029",x"c0e00015",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e007ff",x"f0800002",x"b0000000",
		x"c0e00055",x"c1800cff",x"c1a015ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28dffff",x"f14001ff",x"b0000000",
		x"c0e00035",x"c18002ff",x"c1a00dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2afffff",x"f14003ff",x"b0000000",
		x"c0e00075",x"c1800aff",x"c1a01dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2bfffff",x"f12001bf",x"b0000000",
		x"400000dc",x"c0e00009",x"c0e00049",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e013ff",x"f0a00004",x"b0000000",
		x"400000dd",x"c1000011",x"c1000091",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20023ff",x"f0c00008",x"b0000000",
		x"400000de",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200041",x"f1000020",x"b0000000",
		x"c120001f",x"c14001df",x"c14003df",x"c1a005ff",x"c1a015ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c01fff",x"f10000bf",x"b0000000",
		x"c120011f",x"c140003f",x"c140023f",x"c1a00dff",x"c1a01dff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e03fff",x"f100007f",x"b0000000",
		x"c120009f",x"c140013f",x"c140033f",x"c1a003ff",x"c1a013ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e07fff",x"f10000ff",x"b0000000",
		x"c0c00013",x"c100004f",x"c10000cf",x"c18006ff",x"c1800eff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c02fff",x"f0e0005f",x"b0000000",
		x"c0c00033",x"c100002f",x"c10000af",x"c18001ff",x"c18009ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c01fff",x"f0e0003f",x"b0000000",
		x"400000df",x"c0a00009",x"c0a00019",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c160037f",x"f080000d",x"b0000000",
		x"c0a00005",x"c10000f7",x"c100000f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a01bff",x"f0e0002f",x"b0000000",
		x"c0a00015",x"c100008f",x"c100004f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c007ff",x"f100001f",x"b0000000",
		x"c0a0000d",x"c10000cf",x"c100002f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c027ff",x"f0e0006f",x"b0000000",
		x"c10000af",x"c160077f",x"c16000ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200ffff",x"f14003ff",x"b0000000",
		x"400000e0",x"c0a00009",x"c0a00019",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18001ff",x"f0800009",x"b0000000",
		x"c0a00005",x"c120012f",x"c12000af",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e077ff",x"f0e00037",x"b0000000",
		x"c0a00015",x"c12001af",x"c120006f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e00fff",x"f0e00077",x"b0000000",
		x"c0a0000d",x"c120016f",x"c12000ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e04fff",x"f0e0000f",x"b0000000",
		x"400000e1",x"c0a00013",x"400000e2",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a01bff",x"f0600005",x"b0000000",
		x"400000e3",x"c14003ef",x"c140001f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220dfff",x"f100006f",x"b0000000",
		x"400000e4",x"400000e5",x"c0c00039",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c027ff",x"f080000a",x"b0000000",
		x"400000e6",x"c160023f",x"c160063f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28f7fff",x"f14003df",x"b0000000",
		x"400000e7",x"c160013f",x"c160053f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c280ffff",x"f140003f",x"b0000000",
		x"400000e8",x"c160033f",x"c160073f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c288ffff",x"f140023f",x"b0000000",
		x"400000e9",x"c16000bf",x"c16004bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c284ffff",x"f140013f",x"b0000000",
		x"400000ea",x"c0c00019",x"c0e0000d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e047ff",x"f0a0000a",x"b0000000",
		x"400000eb",x"c0e00029",x"c0e00069",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e053ff",x"f0a00014",x"b0000000",
		x"400000ec",x"c1000051",x"c10000d1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200a3ff",x"f0c00028",x"b0000000",
		x"400000ed",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200141",x"f10000a0",x"b0000000",
		x"400000ee",x"c0a0001d",x"400000ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16004ff",x"f0a00003",x"b0000000",
		x"400000f0",x"c0a0001d",x"400000f1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18009ff",x"f0800005",x"b0000000",
		x"400000f2",x"c0a0000b",x"400000f3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a007ff",x"f0800003",x"b0000000",
		x"400000f4",x"c140021f",x"c140011f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c241dfff",x"f12000ef",x"b0000000",
		x"400000f5",x"c140031f",x"c140009f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c243dfff",x"f12001ef",x"b0000000",
		x"400000f6",x"400000f7",x"c0c00005",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c017ff",x"f0800006",x"b0000000",
		x"400000f8",x"c16002bf",x"c16006bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28cffff",x"f140033f",x"b0000000",
		x"c0c00025",x"c16001bf",x"c16005bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c282ffff",x"f14000bf",x"b0000000",
		x"c0c00015",x"c16003bf",x"c16007bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28affff",x"f14002bf",x"b0000000",
		x"c0c00035",x"c160007f",x"c160047f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c286ffff",x"f14001bf",x"b0000000",
		x"400000f9",x"c160027f",x"c160067f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28effff",x"f14003bf",x"b0000000",
		x"400000fa",x"c0c00039",x"c0e0004d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e027ff",x"f0a0001a",x"b0000000",
		x"400000fb",x"c0e00019",x"c0e00059",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e033ff",x"f0a0000c",x"b0000000",
		x"400000fc",x"c1000031",x"c10000b1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20063ff",x"f0c00018",x"b0000000",
		x"400000fd",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000c1",x"f1000060",x"b0000000",
		x"400000fe",x"400000ff",x"40000100",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16002ff",x"f0a00013",x"b0000000",
		x"40000101",x"c12000ef",x"c12001ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c017ff",x"f100009f",x"b0000000",
		x"40000102",x"c0a00003",x"40000103",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18005ff",x"f080000d",x"b0000000",
		x"40000104",x"c12001ef",x"c140025f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2006fff",x"f10000af",x"b0000000",
		x"40000105",x"40000106",x"40000107",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a017ff",x"f080000b",x"b0000000",
		x"40000108",x"c140029f",x"c160007f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2403fff",x"f120001f",x"b0000000",
		x"40000109",x"c140019f",x"c160047f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2423fff",x"f120011f",x"b0000000",
		x"4000010a",x"c140039f",x"c160027f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2413fff",x"f120009f",x"b0000000",
		x"4000010b",x"c0c0000d",x"c0c0002d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e037ff",x"f080000e",x"b0000000",
		x"c0c0001d",x"c160017f",x"c160057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c281ffff",x"f140007f",x"b0000000",
		x"c0c0003d",x"c160037f",x"c160077f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c289ffff",x"f140027f",x"b0000000",
		x"c0c00003",x"c16000ff",x"c18004ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c285ffff",x"f140017f",x"b0000000",
		x"4000010c",x"c0c00005",x"c0e0002d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e067ff",x"f0a00006",x"b0000000",
		x"4000010d",x"c0e00039",x"c0e00079",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e073ff",x"f0a0001c",x"b0000000",
		x"4000010e",x"c1000071",x"c10000f1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200e3ff",x"f0c00038",x"b0000000",
		x"4000010f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001c1",x"f10000e0",x"b0000000",
		x"40000110",x"c0c00003",x"c0c00023",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c16006ff",x"f0a0000b",x"b0000000",
		x"40000111",x"c120001f",x"c120011f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c037ff",x"f100005f",x"b0000000",
		x"c0c00013",x"c120009f",x"c120019f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e06fff",x"f10000df",x"b0000000",
		x"c0c00033",x"c120005f",x"c120015f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1c00fff",x"f100003f",x"b0000000",
		x"40000112",x"40000113",x"40000114",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800dff",x"f0800003",x"b0000000",
		x"40000115",x"c120001f",x"c140015f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200efff",x"f100006f",x"b0000000",
		x"40000116",x"c120011f",x"c140035f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2001fff",x"f10000ef",x"b0000000",
		x"c0200000",x"40000117",x"40000118",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1a00fff",x"f0800007",x"b0000000",
		x"40000119",x"c140005f",x"c140025f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2433fff",x"f120019f",x"b0000000",
		x"4000011a",x"c140015f",x"c160067f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c240bfff",x"f120005f",x"b0000000",
		x"c0c0001b",x"c140035f",x"c160017f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c242bfff",x"f120015f",x"b0000000",
		x"c0c0003b",x"c14000df",x"c160057f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c241bfff",x"f12000df",x"b0000000",
		x"c0c00007",x"c14002df",x"c160037f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c243bfff",x"f12001df",x"b0000000",
		x"4000011b",x"c0c00023",x"c0c00013",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e077ff",x"f0800001",x"b0000000",
		x"4000011c",x"c0c00025",x"c0e0006d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e017ff",x"f0a00016",x"b0000000",
		x"4000011d",x"c0e00005",x"c0e00045",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e00bff",x"f0a00002",x"b0000000",
		x"4000011e",x"c1000009",x"c1000089",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20013ff",x"f0c00004",x"b0000000",
		x"4000011f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200021",x"f1000010",x"b0000000",
		x"c0600000",x"c0c0000b",x"40000120",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800dff",x"f0a0001b",x"b0000000",
		x"c0c0002b",x"c12000df",x"c12001df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e01fff",x"f10000bf",x"b0000000",
		x"40000121",x"40000122",x"c0c00013",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c18003ff",x"f0a0000b",x"b0000000",
		x"40000123",x"c120009f",x"c14000df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2009fff",x"f100001f",x"b0000000",
		x"c0c00033",x"c14002df",x"c14001df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2207fff",x"f100009f",x"b0000000",
		x"c0c0000b",x"c14003df",x"c140003f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2005fff",x"f100005f",x"b0000000",
		x"c0c0002b",x"c140023f",x"c140013f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200dfff",x"f10000df",x"b0000000",
		x"40000124",x"c14001df",x"c14003df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2407fff",x"f120003f",x"b0000000",
		x"c0c00027",x"c140003f",x"c160077f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2427fff",x"f120013f",x"b0000000",
		x"40000125",x"c140023f",x"c140013f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2417fff",x"f12000bf",x"b0000000",
		x"c0c00017",x"c140033f",x"c16000ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2437fff",x"f12001bf",x"b0000000",
		x"40000126",x"c0c00033",x"c0c0000b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e00fff",x"f0800009",x"b0000000",
		x"40000127",x"40000128",x"c0e0001d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e057ff",x"f0a0000e",x"b0000000",
		x"40000129",x"c0e00025",x"c1000013",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e04bff",x"f0a00012",x"b0000000",
		x"4000012a",x"c1000049",x"c10000c9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20093ff",x"f0c00024",x"b0000000",
		x"4000012b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200121",x"f1000090",x"b0000000",
		x"4000012c",x"c14003bf",x"c140007f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e05fff",x"f120017f",x"b0000000",
		x"c0400000",x"4000012d",x"c0c0001b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1800bff",x"f0a0001b",x"b0000000",
		x"4000012e",x"c140033f",x"c14000bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2003fff",x"f100003f",x"b0000000",
		x"4000012f",x"c120019f",x"c14002bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200bfff",x"f10000bf",x"b0000000",
		x"40000130",x"c14000bf",x"c16004ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c240ffff",x"f120007f",x"b0000000",
		x"40000131",x"c14002bf",x"c16002ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c242ffff",x"f120017f",x"b0000000",
		x"40000132",x"c0c0002b",x"c0c0001b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e04fff",x"f0800005",x"b0000000",
		x"40000133",x"40000134",x"c0e0005d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e037ff",x"f0a0001e",x"b0000000",
		x"40000135",x"c18006ff",x"c1a003ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c283ffff",x"f120007f",x"b0000000",
		x"40000136",x"c0e00065",x"c1000093",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e02bff",x"f0a0000a",x"b0000000",
		x"40000137",x"c1000029",x"c10000a9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20053ff",x"f0c00014",x"b0000000",
		x"40000138",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000a1",x"f1000050",x"b0000000",
		x"c0e00037",x"c140027f",x"c140017f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e03fff",x"f12000ff",x"b0000000",
		x"c0c0003b",x"c14001bf",x"c14003bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2217fff",x"f12000ff",x"b0000000",
		x"c0c00007",x"c140007f",x"c140027f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220ffff",x"f12001ff",x"b0000000",
		x"c0c00027",x"c140017f",x"c140037f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221ffff",x"f100007f",x"b0000000",
		x"c0c00037",x"c14001bf",x"c16006ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c241ffff",x"f12000ff",x"b0000000",
		x"c0c0000f",x"c14003bf",x"c16001ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c243ffff",x"f12001ff",x"b0000000",
		x"40000139",x"c0c0003b",x"4000013a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e02fff",x"f080000d",x"b0000000",
		x"4000013b",x"c0e0003d",x"c0e0007d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e077ff",x"f0a00001",x"b0000000",
		x"c0e00003",x"c1800eff",x"c1a013ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28bffff",x"f120017f",x"b0000000",
		x"c0e00043",x"c18001ff",x"c1a00bff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c287ffff",x"f12000ff",x"b0000000",
		x"4000013c",x"c0e00015",x"c1000053",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e06bff",x"f0a0001a",x"b0000000",
		x"4000013d",x"c1000069",x"c10000e9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200d3ff",x"f0c00034",x"b0000000",
		x"4000013e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001a1",x"f10000d0",x"b0000000",
		x"4000013f",x"c0c00007",x"40000140",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e06fff",x"f0800003",x"b0000000",
		x"40000141",x"c1800cff",x"c18002ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28dffff",x"f140037f",x"b0000000",
		x"40000142",x"c0e00023",x"c0e00063",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e00fff",x"f0a00011",x"b0000000",
		x"40000143",x"c0e00055",x"c10000d3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e01bff",x"f0a00006",x"b0000000",
		x"40000144",x"c1000019",x"c1000099",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20033ff",x"f0c0000c",x"b0000000",
		x"40000145",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200061",x"f1000030",x"b0000000",
		x"40000146",x"c0c00027",x"40000147",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e01fff",x"f080000b",x"b0000000",
		x"c0e0000f",x"c1800aff",x"c18006ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c283ffff",x"f14000ff",x"b0000000",
		x"40000148",x"c1800eff",x"c18001ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28bffff",x"f14002ff",x"b0000000",
		x"40000149",x"c0e00013",x"c0e00053",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2004fff",x"f0a00009",x"b0000000",
		x"4000014a",x"c0e00035",x"c1000033",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e05bff",x"f0a00016",x"b0000000",
		x"4000014b",x"c1000059",x"c10000d9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200b3ff",x"f0c0002c",x"b0000000",
		x"4000014c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200161",x"f10000b0",x"b0000000",
		x"4000014d",x"c0c00017",x"c0e0004f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e05fff",x"f0800007",x"b0000000",
		x"c0e0002f",x"c18009ff",x"c18005ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c287ffff",x"f14001ff",x"b0000000",
		x"c0e0006f",x"c1800dff",x"c18003ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c28fffff",x"f14003ff",x"b0000000",
		x"4000014e",x"c0e00033",x"c0e00073",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200cfff",x"f0a00019",x"b0000000",
		x"4000014f",x"c0e00075",x"c10000b3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e03bff",x"f0a0000e",x"b0000000",
		x"40000150",x"c1000039",x"c10000b9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20073ff",x"f0c0001c",x"b0000000",
		x"40000151",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000e1",x"f1000070",x"b0000000",
		x"c0200000",x"c0c00037",x"c0e0001f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e03fff",x"f0a0000f",x"b0000000",
		x"40000152",x"c0e0000b",x"c0e0004b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2002fff",x"f0a00005",x"b0000000",
		x"40000153",x"c0e0000d",x"c1000073",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e07bff",x"f0a0001e",x"b0000000",
		x"40000154",x"c1000079",x"c10000f9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200f3ff",x"f0c0003c",x"b0000000",
		x"40000155",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001e1",x"f10000f0",x"b0000000",
		x"40000156",x"c0e0002b",x"c0e0006b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200afff",x"f0a00015",x"b0000000",
		x"40000157",x"c0e0004d",x"c10000f3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e007ff",x"f0a00001",x"b0000000",
		x"40000158",x"c1000005",x"c1000085",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2000bff",x"f0c00002",x"b0000000",
		x"40000159",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200011",x"f1000008",x"b0000000",
		x"4000015a",x"c0e0001b",x"c0e0005b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2006fff",x"f0a0000d",x"b0000000",
		x"4000015b",x"c0e0002d",x"c100000b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1e047ff",x"f0a00011",x"b0000000",
		x"4000015c",x"c1000045",x"c10000c5",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2008bff",x"f0c00022",x"b0000000",
		x"4000015d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200111",x"f1000088",x"b0000000",
		x"4000015e",x"c0e0003b",x"c0e0007b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200efff",x"f0a0001d",x"b0000000",
		x"4000015f",x"c0e0006d",x"c100008b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20027ff",x"f0c00009",x"b0000000",
		x"40000160",x"c1000025",x"c10000a5",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2004bff",x"f0c00012",x"b0000000",
		x"40000161",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200091",x"f1000048",x"b0000000",
		x"40000162",x"c0e00007",x"c0e00047",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2001fff",x"f0a00003",x"b0000000",
		x"40000163",x"c0e0001d",x"c100004b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200a7ff",x"f0c00029",x"b0000000",
		x"40000164",x"c1000065",x"c10000e5",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200cbff",x"f0c00032",x"b0000000",
		x"40000165",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200191",x"f10000c8",x"b0000000",
		x"40000166",x"c0e00027",x"c0e00067",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2009fff",x"f0a00013",x"b0000000",
		x"40000167",x"c0e0005d",x"c10000cb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20067ff",x"f0c00019",x"b0000000",
		x"40000168",x"c1000015",x"c1000095",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2002bff",x"f0c0000a",x"b0000000",
		x"40000169",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200051",x"f1000028",x"b0000000",
		x"4000016a",x"c0e00017",x"c0e00057",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2005fff",x"f0a0000b",x"b0000000",
		x"4000016b",x"c0e0003d",x"c100002b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200e7ff",x"f0c00039",x"b0000000",
		x"4000016c",x"c1000055",x"c120006b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200abff",x"f0c0002a",x"b0000000",
		x"4000016d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200151",x"f10000a8",x"b0000000",
		x"4000016e",x"c0e00037",x"c0e00077",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200dfff",x"f0a0001b",x"b0000000",
		x"4000016f",x"c0e0007d",x"c10000ab",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20017ff",x"f0c00005",x"b0000000",
		x"40000170",x"c10000d5",x"c120016b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2006bff",x"f0c0001a",x"b0000000",
		x"40000171",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000d1",x"f1000068",x"b0000000",
		x"40000172",x"c0e0000f",x"c0e0004f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2003fff",x"f0a00007",x"b0000000",
		x"40000173",x"c0e00003",x"c100006b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20097ff",x"f0c00025",x"b0000000",
		x"40000174",x"c1000035",x"c12000eb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200ebff",x"f0c0003a",x"b0000000",
		x"40000175",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001d1",x"f10000e8",x"b0000000",
		x"40000176",x"c0e0002f",x"c0e0006f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200bfff",x"f0a00017",x"b0000000",
		x"40000177",x"c0e00043",x"c10000eb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20057ff",x"f0c00015",x"b0000000",
		x"40000178",x"c10000b5",x"c12001eb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2001bff",x"f0c00006",x"b0000000",
		x"40000179",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200031",x"f1000018",x"b0000000",
		x"4000017a",x"c0e0001f",x"c0e0005f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2007fff",x"f0a0000f",x"b0000000",
		x"4000017b",x"c0e00023",x"c100001b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200d7ff",x"f0c00035",x"b0000000",
		x"4000017c",x"c1000075",x"c120001b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2009bff",x"f0c00026",x"b0000000",
		x"4000017d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200131",x"f1000098",x"b0000000",
		x"c0200000",x"c0e0003f",x"c100007f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220ffff",x"f0c0001f",x"b0000000",
		x"4000017e",x"c0e00063",x"c100009b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20037ff",x"f0c0000d",x"b0000000",
		x"4000017f",x"c10000f5",x"c120011b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2005bff",x"f0c00016",x"b0000000",
		x"40000180",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000b1",x"f1000058",x"b0000000",
		x"40000181",x"c100005b",x"c10000db",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200b7ff",x"f0c0002d",x"b0000000",
		x"40000182",x"c100000d",x"c120009b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200dbff",x"f0c00036",x"b0000000",
		x"40000183",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001b1",x"f10000d8",x"b0000000",
		x"40000184",x"c100003b",x"c10000bb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20077ff",x"f0c0001d",x"b0000000",
		x"40000185",x"c100008d",x"c120019b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2003bff",x"f0c0000e",x"b0000000",
		x"40000186",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200071",x"f1000038",x"b0000000",
		x"40000187",x"c100007b",x"c10000fb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200f7ff",x"f0c0003d",x"b0000000",
		x"40000188",x"c100004d",x"c120005b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200bbff",x"f0c0002e",x"b0000000",
		x"40000189",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200171",x"f10000b8",x"b0000000",
		x"4000018a",x"c1000007",x"c1000087",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2000fff",x"f0c00003",x"b0000000",
		x"4000018b",x"c10000cd",x"c120015b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2007bff",x"f0c0001e",x"b0000000",
		x"4000018c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000f1",x"f1000078",x"b0000000",
		x"4000018d",x"c1000047",x"c10000c7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2008fff",x"f0c00023",x"b0000000",
		x"4000018e",x"c100002d",x"c12000db",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200fbff",x"f0c0003e",x"b0000000",
		x"4000018f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001f1",x"f10000f8",x"b0000000",
		x"40000190",x"c1000027",x"c10000a7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2004fff",x"f0c00013",x"b0000000",
		x"40000191",x"c10000ad",x"c12001db",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20007ff",x"f0c00001",x"b0000000",
		x"40000192",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200009",x"f1000004",x"b0000000",
		x"40000193",x"c1000067",x"c10000e7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200cfff",x"f0c00033",x"b0000000",
		x"40000194",x"c100006d",x"c120003b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20087ff",x"f0c00021",x"b0000000",
		x"40000195",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200109",x"f1000084",x"b0000000",
		x"40000196",x"c1000017",x"c1000097",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2002fff",x"f0c0000b",x"b0000000",
		x"40000197",x"c10000ed",x"c120013b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20047ff",x"f0c00011",x"b0000000",
		x"40000198",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200089",x"f1000044",x"b0000000",
		x"40000199",x"c1000057",x"c10000d7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200afff",x"f0c0002b",x"b0000000",
		x"4000019a",x"c100001d",x"c12000bb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200c7ff",x"f0c00031",x"b0000000",
		x"4000019b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200189",x"f10000c4",x"b0000000",
		x"4000019c",x"c1000037",x"c10000b7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2006fff",x"f0c0001b",x"b0000000",
		x"4000019d",x"c100009d",x"c12001bb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20027ff",x"f0c00009",x"b0000000",
		x"4000019e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200049",x"f1000024",x"b0000000",
		x"4000019f",x"c1000077",x"c10000f7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200efff",x"f0c0003b",x"b0000000",
		x"400001a0",x"c100005d",x"c120007b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200a7ff",x"f0c00029",x"b0000000",
		x"400001a1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200149",x"f10000a4",x"b0000000",
		x"400001a2",x"c100000f",x"c100008f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2001fff",x"f0c00007",x"b0000000",
		x"400001a3",x"c10000dd",x"c120017b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20067ff",x"f0c00019",x"b0000000",
		x"400001a4",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000c9",x"f1000064",x"b0000000",
		x"400001a5",x"c100004f",x"c10000cf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2009fff",x"f0c00027",x"b0000000",
		x"400001a6",x"c100003d",x"c12000fb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200e7ff",x"f0c00039",x"b0000000",
		x"400001a7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001c9",x"f10000e4",x"b0000000",
		x"400001a8",x"c100002f",x"c10000af",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2005fff",x"f0c00017",x"b0000000",
		x"400001a9",x"c10000bd",x"c12001fb",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20017ff",x"f0c00005",x"b0000000",
		x"400001aa",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200029",x"f1000014",x"b0000000",
		x"400001ab",x"c100006f",x"c10000ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200dfff",x"f0c00037",x"b0000000",
		x"400001ac",x"c100007d",x"c1200007",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20097ff",x"f0c00025",x"b0000000",
		x"400001ad",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200129",x"f1000094",x"b0000000",
		x"400001ae",x"c100001f",x"c100009f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2003fff",x"f0c0000f",x"b0000000",
		x"400001af",x"c10000fd",x"c1200107",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c20057ff",x"f0c00015",x"b0000000",
		x"400001b0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000a9",x"f1000054",x"b0000000",
		x"400001b1",x"c100005f",x"c10000df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c200bfff",x"f0c0002f",x"b0000000",
		x"400001b2",x"c1000003",x"c1200087",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220d7ff",x"f0e00035",x"b0000000",
		x"400001b3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001a9",x"f10000d4",x"b0000000",
		x"400001b4",x"c100003f",x"c10000bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2007fff",x"f0c0001f",x"b0000000",
		x"400001b5",x"c1000083",x"c1200187",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221d7ff",x"f0e00075",x"b0000000",
		x"400001b6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200069",x"f1000034",x"b0000000",
		x"c0200000",x"c100007f",x"c12000ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220ffff",x"f0e0003f",x"b0000000",
		x"400001b7",x"c1000043",x"c1200047",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c22037ff",x"f0e0000d",x"b0000000",
		x"400001b8",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200169",x"f10000b4",x"b0000000",
		x"400001b9",x"c10000c3",x"c1200147",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c22137ff",x"f0e0004d",x"b0000000",
		x"400001ba",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000e9",x"f1000074",x"b0000000",
		x"400001bb",x"c1000023",x"c12000c7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220b7ff",x"f0e0002d",x"b0000000",
		x"400001bc",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001e9",x"f10000f4",x"b0000000",
		x"400001bd",x"c10000a3",x"c12001c7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221b7ff",x"f0e0006d",x"b0000000",
		x"400001be",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200019",x"f100000c",x"b0000000",
		x"400001bf",x"c1000063",x"c1200027",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c22077ff",x"f0e0001d",x"b0000000",
		x"400001c0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200119",x"f100008c",x"b0000000",
		x"400001c1",x"c10000e3",x"c1200127",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c22177ff",x"f0e0005d",x"b0000000",
		x"400001c2",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200099",x"f100004c",x"b0000000",
		x"400001c3",x"c1000013",x"c12000a7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220f7ff",x"f0e0003d",x"b0000000",
		x"400001c4",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200199",x"f10000cc",x"b0000000",
		x"400001c5",x"c1000093",x"c12001a7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221f7ff",x"f0e0007d",x"b0000000",
		x"400001c6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200059",x"f100002c",x"b0000000",
		x"400001c7",x"c1000053",x"c1200067",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2200fff",x"f0e00003",x"b0000000",
		x"400001c8",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200159",x"f10000ac",x"b0000000",
		x"400001c9",x"c10000d3",x"c1200167",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2210fff",x"f0e00043",x"b0000000",
		x"400001ca",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000d9",x"f100006c",x"b0000000",
		x"400001cb",x"c1000033",x"c12000e7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2208fff",x"f0e00023",x"b0000000",
		x"400001cc",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001d9",x"f10000ec",x"b0000000",
		x"400001cd",x"c10000b3",x"c12001e7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2218fff",x"f0e00063",x"b0000000",
		x"400001ce",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200039",x"f100001c",x"b0000000",
		x"400001cf",x"c1000073",x"c1200017",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2204fff",x"f0e00013",x"b0000000",
		x"400001d0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200139",x"f100009c",x"b0000000",
		x"400001d1",x"c10000f3",x"c1200117",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2214fff",x"f0e00053",x"b0000000",
		x"400001d2",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000b9",x"f100005c",x"b0000000",
		x"400001d3",x"c100000b",x"c1200097",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220cfff",x"f0e00033",x"b0000000",
		x"400001d4",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001b9",x"f10000dc",x"b0000000",
		x"400001d5",x"c100008b",x"c1200197",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221cfff",x"f0e00073",x"b0000000",
		x"400001d6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200079",x"f100003c",x"b0000000",
		x"400001d7",x"c100004b",x"c1200057",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2202fff",x"f0e0000b",x"b0000000",
		x"400001d8",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200179",x"f10000bc",x"b0000000",
		x"400001d9",x"c10000cb",x"c1200157",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2212fff",x"f0e0004b",x"b0000000",
		x"400001da",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000f9",x"f100007c",x"b0000000",
		x"400001db",x"c100002b",x"c12000d7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220afff",x"f0e0002b",x"b0000000",
		x"400001dc",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001f9",x"f10000fc",x"b0000000",
		x"400001dd",x"c10000ab",x"c12001d7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221afff",x"f0e0006b",x"b0000000",
		x"400001de",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200005",x"f1000002",x"b0000000",
		x"400001df",x"c1200037",x"c1200137",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2206fff",x"f0e0001b",x"b0000000",
		x"400001e0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200105",x"f1000082",x"b0000000",
		x"400001e1",x"c12000b7",x"c12001b7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2216fff",x"f0e0005b",x"b0000000",
		x"400001e2",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200085",x"f1000042",x"b0000000",
		x"400001e3",x"c1200077",x"c1200177",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220efff",x"f0e0003b",x"b0000000",
		x"400001e4",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200185",x"f10000c2",x"b0000000",
		x"400001e5",x"c12000f7",x"c12001f7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221efff",x"f0e0007b",x"b0000000",
		x"400001e6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200045",x"f1000022",x"b0000000",
		x"400001e7",x"c120000f",x"c120010f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2201fff",x"f0e00007",x"b0000000",
		x"400001e8",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200145",x"f10000a2",x"b0000000",
		x"400001e9",x"c120008f",x"c120018f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2211fff",x"f0e00047",x"b0000000",
		x"400001ea",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000c5",x"f1000062",x"b0000000",
		x"400001eb",x"c120004f",x"c120014f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2209fff",x"f0e00027",x"b0000000",
		x"400001ec",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001c5",x"f10000e2",x"b0000000",
		x"400001ed",x"c12000cf",x"c12001cf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2219fff",x"f0e00067",x"b0000000",
		x"400001ee",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200025",x"f1000012",x"b0000000",
		x"400001ef",x"c120002f",x"c120012f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2205fff",x"f0e00017",x"b0000000",
		x"400001f0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200125",x"f1000092",x"b0000000",
		x"400001f1",x"c12000af",x"c12001af",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2215fff",x"f0e00057",x"b0000000",
		x"400001f2",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000a5",x"f1000052",x"b0000000",
		x"400001f3",x"c120006f",x"c120016f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220dfff",x"f0e00037",x"b0000000",
		x"400001f4",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001a5",x"f10000d2",x"b0000000",
		x"400001f5",x"c12000ef",x"c12001ef",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221dfff",x"f0e00077",x"b0000000",
		x"400001f6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200065",x"f1000032",x"b0000000",
		x"400001f7",x"c120001f",x"c120011f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2203fff",x"f0e0000f",x"b0000000",
		x"400001f8",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200165",x"f10000b2",x"b0000000",
		x"400001f9",x"c120009f",x"c120019f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2213fff",x"f0e0004f",x"b0000000",
		x"400001fa",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000e5",x"f1000072",x"b0000000",
		x"400001fb",x"c120005f",x"c120015f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220bfff",x"f0e0002f",x"b0000000",
		x"400001fc",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001e5",x"f10000f2",x"b0000000",
		x"400001fd",x"c12000df",x"c12001df",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221bfff",x"f0e0006f",x"b0000000",
		x"400001fe",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200015",x"f100000a",x"b0000000",
		x"400001ff",x"c120003f",x"c120013f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2207fff",x"f0e0001f",x"b0000000",
		x"40000200",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200115",x"f100008a",x"b0000000",
		x"40000201",x"c12000bf",x"c12001bf",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c2217fff",x"f0e0005f",x"b0000000",
		x"40000202",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200095",x"f100004a",x"b0000000",
		x"40000203",x"c120007f",x"c120017f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c220ffff",x"f0e0003f",x"b0000000",
		x"40000204",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200195",x"f10000ca",x"b0000000",
		x"c0200000",x"c12000ff",x"c14001ff",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c221ffff",x"f0e0007f",x"b0000000",
		x"40000205",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200055",x"f100002a",x"b0000000",
		x"40000206",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200155",x"f10000aa",x"b0000000",
		x"40000207",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000d5",x"f100006a",x"b0000000",
		x"40000208",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001d5",x"f10000ea",x"b0000000",
		x"40000209",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200035",x"f100001a",x"b0000000",
		x"4000020a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200135",x"f100009a",x"b0000000",
		x"4000020b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000b5",x"f100005a",x"b0000000",
		x"4000020c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001b5",x"f10000da",x"b0000000",
		x"4000020d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200075",x"f100003a",x"b0000000",
		x"4000020e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200175",x"f10000ba",x"b0000000",
		x"4000020f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000f5",x"f100007a",x"b0000000",
		x"40000210",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001f5",x"f10000fa",x"b0000000",
		x"40000211",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120000d",x"f1000006",x"b0000000",
		x"40000212",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120010d",x"f1000086",x"b0000000",
		x"40000213",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120008d",x"f1000046",x"b0000000",
		x"40000214",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120018d",x"f10000c6",x"b0000000",
		x"40000215",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120004d",x"f1000026",x"b0000000",
		x"40000216",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120014d",x"f10000a6",x"b0000000",
		x"40000217",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000cd",x"f1000066",x"b0000000",
		x"40000218",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001cd",x"f10000e6",x"b0000000",
		x"40000219",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120002d",x"f1000016",x"b0000000",
		x"4000021a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120012d",x"f1000096",x"b0000000",
		x"4000021b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000ad",x"f1000056",x"b0000000",
		x"4000021c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001ad",x"f10000d6",x"b0000000",
		x"4000021d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120006d",x"f1000036",x"b0000000",
		x"4000021e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120016d",x"f10000b6",x"b0000000",
		x"4000021f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000ed",x"f1000076",x"b0000000",
		x"40000220",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001ed",x"f10000f6",x"b0000000",
		x"40000221",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120001d",x"f100000e",x"b0000000",
		x"40000222",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120011d",x"f100008e",x"b0000000",
		x"40000223",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120009d",x"f100004e",x"b0000000",
		x"40000224",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120019d",x"f10000ce",x"b0000000",
		x"40000225",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120005d",x"f100002e",x"b0000000",
		x"40000226",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120015d",x"f10000ae",x"b0000000",
		x"40000227",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000dd",x"f100006e",x"b0000000",
		x"40000228",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001dd",x"f10000ee",x"b0000000",
		x"40000229",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120003d",x"f100001e",x"b0000000",
		x"4000022a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120013d",x"f100009e",x"b0000000",
		x"4000022b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000bd",x"f100005e",x"b0000000",
		x"4000022c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001bd",x"f10000de",x"b0000000",
		x"4000022d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120007d",x"f100003e",x"b0000000",
		x"4000022e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120017d",x"f10000be",x"b0000000",
		x"4000022f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000fd",x"f100007e",x"b0000000",
		x"40000230",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001fd",x"f10000fe",x"b0000000",
		x"40000231",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200003",x"f1000001",x"b0000000",
		x"40000232",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200103",x"f1000081",x"b0000000",
		x"40000233",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200083",x"f1000041",x"b0000000",
		x"40000234",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200183",x"f10000c1",x"b0000000",
		x"40000235",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200043",x"f1000021",x"b0000000",
		x"40000236",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200143",x"f10000a1",x"b0000000",
		x"40000237",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000c3",x"f1000061",x"b0000000",
		x"40000238",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001c3",x"f10000e1",x"b0000000",
		x"40000239",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200023",x"f1000011",x"b0000000",
		x"4000023a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200123",x"f1000091",x"b0000000",
		x"4000023b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000a3",x"f1000051",x"b0000000",
		x"4000023c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001a3",x"f10000d1",x"b0000000",
		x"4000023d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200063",x"f1000031",x"b0000000",
		x"4000023e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200163",x"f10000b1",x"b0000000",
		x"4000023f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000e3",x"f1000071",x"b0000000",
		x"40000240",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001e3",x"f10000f1",x"b0000000",
		x"40000241",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200013",x"f1000009",x"b0000000",
		x"40000242",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200113",x"f1000089",x"b0000000",
		x"40000243",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200093",x"f1000049",x"b0000000",
		x"40000244",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200193",x"f10000c9",x"b0000000",
		x"40000245",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200053",x"f1000029",x"b0000000",
		x"40000246",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200153",x"f10000a9",x"b0000000",
		x"40000247",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000d3",x"f1000069",x"b0000000",
		x"40000248",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001d3",x"f10000e9",x"b0000000",
		x"40000249",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200033",x"f1000019",x"b0000000",
		x"4000024a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200133",x"f1000099",x"b0000000",
		x"4000024b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000b3",x"f1000059",x"b0000000",
		x"4000024c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001b3",x"f10000d9",x"b0000000",
		x"4000024d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200073",x"f1000039",x"b0000000",
		x"4000024e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200173",x"f10000b9",x"b0000000",
		x"4000024f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000f3",x"f1000079",x"b0000000",
		x"40000250",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001f3",x"f10000f9",x"b0000000",
		x"40000251",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120000b",x"f1000005",x"b0000000",
		x"40000252",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120010b",x"f1000085",x"b0000000",
		x"40000253",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120008b",x"f1000045",x"b0000000",
		x"40000254",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120018b",x"f10000c5",x"b0000000",
		x"40000255",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120004b",x"f1000025",x"b0000000",
		x"40000256",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120014b",x"f10000a5",x"b0000000",
		x"40000257",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000cb",x"f1000065",x"b0000000",
		x"40000258",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001cb",x"f10000e5",x"b0000000",
		x"40000259",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120002b",x"f1000015",x"b0000000",
		x"4000025a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120012b",x"f1000095",x"b0000000",
		x"4000025b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000ab",x"f1000055",x"b0000000",
		x"4000025c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001ab",x"f10000d5",x"b0000000",
		x"4000025d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120006b",x"f1000035",x"b0000000",
		x"4000025e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120016b",x"f10000b5",x"b0000000",
		x"4000025f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000eb",x"f1000075",x"b0000000",
		x"40000260",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001eb",x"f10000f5",x"b0000000",
		x"40000261",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120001b",x"f100000d",x"b0000000",
		x"40000262",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120011b",x"f100008d",x"b0000000",
		x"40000263",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120009b",x"f100004d",x"b0000000",
		x"40000264",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120019b",x"f10000cd",x"b0000000",
		x"40000265",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120005b",x"f100002d",x"b0000000",
		x"40000266",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120015b",x"f10000ad",x"b0000000",
		x"40000267",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000db",x"f100006d",x"b0000000",
		x"40000268",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001db",x"f10000ed",x"b0000000",
		x"40000269",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120003b",x"f100001d",x"b0000000",
		x"4000026a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120013b",x"f100009d",x"b0000000",
		x"4000026b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000bb",x"f100005d",x"b0000000",
		x"4000026c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001bb",x"f10000dd",x"b0000000",
		x"4000026d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120007b",x"f100003d",x"b0000000",
		x"4000026e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120017b",x"f10000bd",x"b0000000",
		x"4000026f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000fb",x"f100007d",x"b0000000",
		x"40000270",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001fb",x"f10000fd",x"b0000000",
		x"40000271",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200007",x"f1000003",x"b0000000",
		x"40000272",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200107",x"f1000083",x"b0000000",
		x"40000273",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200087",x"f1000043",x"b0000000",
		x"40000274",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200187",x"f10000c3",x"b0000000",
		x"40000275",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200047",x"f1000023",x"b0000000",
		x"40000276",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200147",x"f10000a3",x"b0000000",
		x"40000277",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000c7",x"f1000063",x"b0000000",
		x"40000278",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001c7",x"f10000e3",x"b0000000",
		x"40000279",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200027",x"f1000013",x"b0000000",
		x"4000027a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200127",x"f1000093",x"b0000000",
		x"4000027b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000a7",x"f1000053",x"b0000000",
		x"4000027c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001a7",x"f10000d3",x"b0000000",
		x"4000027d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200067",x"f1000033",x"b0000000",
		x"4000027e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200167",x"f10000b3",x"b0000000",
		x"4000027f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000e7",x"f1000073",x"b0000000",
		x"40000280",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001e7",x"f10000f3",x"b0000000",
		x"40000281",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200017",x"f100000b",x"b0000000",
		x"40000282",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200117",x"f100008b",x"b0000000",
		x"40000283",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200097",x"f100004b",x"b0000000",
		x"40000284",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200197",x"f10000cb",x"b0000000",
		x"40000285",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200057",x"f100002b",x"b0000000",
		x"40000286",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200157",x"f10000ab",x"b0000000",
		x"40000287",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000d7",x"f100006b",x"b0000000",
		x"40000288",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001d7",x"f10000eb",x"b0000000",
		x"40000289",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200037",x"f100001b",x"b0000000",
		x"4000028a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200137",x"f100009b",x"b0000000",
		x"4000028b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000b7",x"f100005b",x"b0000000",
		x"4000028c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001b7",x"f10000db",x"b0000000",
		x"4000028d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200077",x"f100003b",x"b0000000",
		x"4000028e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c1200177",x"f10000bb",x"b0000000",
		x"4000028f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000f7",x"f100007b",x"b0000000",
		x"40000290",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001f7",x"f10000fb",x"b0000000",
		x"40000291",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120000f",x"f1000007",x"b0000000",
		x"40000292",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120010f",x"f1000087",x"b0000000",
		x"40000293",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120008f",x"f1000047",x"b0000000",
		x"40000294",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120018f",x"f10000c7",x"b0000000",
		x"40000295",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120004f",x"f1000027",x"b0000000",
		x"40000296",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120014f",x"f10000a7",x"b0000000",
		x"40000297",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000cf",x"f1000067",x"b0000000",
		x"40000298",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001cf",x"f10000e7",x"b0000000",
		x"40000299",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120002f",x"f1000017",x"b0000000",
		x"4000029a",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120012f",x"f1000097",x"b0000000",
		x"4000029b",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000af",x"f1000057",x"b0000000",
		x"4000029c",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001af",x"f10000d7",x"b0000000",
		x"4000029d",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120006f",x"f1000037",x"b0000000",
		x"4000029e",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120016f",x"f10000b7",x"b0000000",
		x"4000029f",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000ef",x"f1000077",x"b0000000",
		x"400002a0",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001ef",x"f10000f7",x"b0000000",
		x"400002a1",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120001f",x"f100000f",x"b0000000",
		x"400002a2",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120011f",x"f100008f",x"b0000000",
		x"400002a3",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120009f",x"f100004f",x"b0000000",
		x"400002a4",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120019f",x"f10000cf",x"b0000000",
		x"400002a5",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120005f",x"f100002f",x"b0000000",
		x"400002a6",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120015f",x"f10000af",x"b0000000",
		x"400002a7",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000df",x"f100006f",x"b0000000",
		x"400002a8",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001df",x"f10000ef",x"b0000000",
		x"400002a9",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120003f",x"f100001f",x"b0000000",
		x"400002aa",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120013f",x"f100009f",x"b0000000",
		x"400002ab",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000bf",x"f100005f",x"b0000000",
		x"400002ac",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001bf",x"f10000df",x"b0000000",
		x"400002ad",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120007f",x"f100003f",x"b0000000",
		x"400002ae",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c120017f",x"f10000bf",x"b0000000",
		x"400002af",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12000ff",x"f100007f",x"b0000000",
		x"c0200000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"b0000000",x"c12001ff",x"f10000ff",x"b0000000"
	);
	
	subtype bin_table_t is std_logic_vector (CONST_LOW_ENTROPY_TABLE_ENTRY_BITS*CONST_INPUT_SYMBOL_AMOUNT-1 downto 0);
    type table_rom_t is array (0 to CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT - 1) of bin_table_t;

    constant CONST_LOW_ENTROPY_CODING_TABLE : table_rom_t := (
		x"f020000040000010c0600000c0600004c060000240000011c0800006c080000e4000001240000013c0a00001c0a00011c0c00005c0c00025c0a00009",
		x"f0200000400000144000001540000016c0600000c0600004c0800002c080000ac0a00006c0a00016c0c0000d40000017b0000000b0000000c0c0002d",
		x"f0200000c04000004000001840000019c0600002c06000064000001a4000001bc0c00019c0c00039b0000000b0000000b0000000b0000000c0c00005",
		x"f02000004000001cc04000004000001d4000001e4000001fc0a0000e40000020b0000000b0000000b0000000b0000000b0000000b0000000c0c00005",
		x"f020000040000021c0400000c0400002c0800001c0800009c0e00013c0e00053b0000000b0000000b0000000b0000000b0000000b0000000c1000027",
		x"f0200000c0200000c040000140000022c0a00003c0a00013b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0e0001b",
		x"f040000040000023400000244000002540000026c0e0000bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120006f",
		x"f02000004000002740000028c060000140000029c12000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c14001bf",
		x"f04000004000002a4000002b4000002cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120006f",
		x"f06000004000002dc0800002c080000ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c140005f",
		x"f06000004000002e4000002fc0a00001b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18005ff",
		x"f080000040000030c0a0000140000031b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c00bff",
		x"f080000040000032c0c00001c0c00021b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e01bff",
		x"f0a000004000003340000034c0e00001b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e003ff",
		x"f0c0000040000035c1000001c1000081b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20003ff",
		x"f100000040000036b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200001",
		x"f0400001c0a000194000003740000038c0c00015c0c00035c0c0000dc0c0002dc0e00013c0e00053c100003bc10000bbc120000fc120010fc100007b",
		x"f0600003c0c0001dc0c0003dc0c00003c0c0002340000039c0e00033c0e00073c10000fbc1000007c120008fc120018fc120004fc120014fc1000087",
		x"f0a00007c0e0000bc0e0004bc0e0002bc1000047c10000c7c1000027c10000a7c12000cfc12001cfc140015fc140035fc160007fc160047fc14000df",
		x"f0a00017c0e0006bc0e0001bc0e0005bc1000067c10000e7c1000017c1000097c120002fc120012fc14002dfc14001dfc160027fc160067fc14003df",
		x"f06000014000003ac0a0000ec0a0001e4000003b4000003cc0c0001dc0c0003dc0e00013c0e00053c12000e7c12001e7b0000000b0000000c100002b",
		x"f0600005c0a00001c0a00011c0a000094000003dc0c000034000003e4000003fc10000abc100006bc1200017c1200117b0000000b0000000c1200097",
		x"f0600003c0a00019c0a00005c0a0001540000040c0c0002340000041c0e00033c10000ebc100001bc1200197c1200057b0000000b0000000c1200157",
		x"f0e0001fc12000d7c12001d7c1200037c14001efc14003efc140001fc140021fc160023fc180017fc1a00dffc1a01dffb0000000b0000000c180097f",
		x"f0600001c080000140000042400000434000004440000045c0e00035c0e00075c100006bc12000f7b0000000b0000000b0000000b0000000c12001f7",
		x"f06000054000004640000047c0a000094000004840000049c0e0000dc0e0004dc10000ebc120000fb0000000b0000000b0000000b0000000c120010f",
		x"f0a00003c0c00025c0e0002dc0e0006dc100001bc100009bc120008fc120018fc16000bfc16004bfb0000000b0000000b0000000b0000000c16002bf",
		x"f0a00013c0e0001dc0e0005dc0e0003dc100005bc10000dbc120004fc120014fc16006bfc16001bfb0000000b0000000b0000000b0000000c16005bf",
		x"f06000014000004ac0800002c080000ac0a0001ec0a00001c0e0002dc0e0006db0000000b0000000b0000000b0000000b0000000b0000000c100006b",
		x"f0600005c08000064000004b4000004c4000004dc0c00025c10000ebc100001bb0000000b0000000b0000000b0000000b0000000b0000000c100009b",
		x"f0800003c0a000114000004e4000004fc0e0001dc0e0005dc1200077c1200177b0000000b0000000b0000000b0000000b0000000b0000000c12000f7",
		x"f0a00007c0a0000940000050c0c00015c0e0003dc0e0007dc12001f7c120000fb0000000b0000000b0000000b0000000b0000000b0000000c14000df",
		x"f0e0000fc0e00003c100005bc10000dbc120010fc120008fc16002bfc16006bfb0000000b0000000b0000000b0000000b0000000b0000000c18002ff",
		x"f04000014000005140000052400000534000005440000055c10000a7c1000067b0000000b0000000b0000000b0000000b0000000b0000000c12000ef",
		x"f0600001400000564000005740000058c0e0005b40000059b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000b7",
		x"f04000024000005ac06000004000005bc0e0004bc0e0002bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120016f",
		x"f0800005c06000044000005cc0a00009c12000efc12001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16001bf",
		x"f080000d4000005dc0a00019c0a00005c120001fc120011fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16005bf",
		x"f100007fc0e0006bc120009fc120019fc1a005ffc1a015ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e03fff",
		x"f0400001c02000004000005e4000005fc12001efc120001fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c160027f",
		x"f08000034000006040000061c0c0000bc160067fc160017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a003ff",
		x"f12000ffc120011fc160057fc160037fc2001fffc220bfffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c241ffff",
		x"f06000024000006240000063c0800004b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120016f",
		x"f0c000074000006440000065c0e0001bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18001ff",
		x"f0c000274000006640000067c0e0005bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18009ff",
		x"f060000440000068c080000640000069b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16000ff",
		x"f06000044000006a4000006bc0a00011b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1800dff",
		x"f100000f4000006cc120002fc14001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2201fff",
		x"f08000084000006d4000006e4000006fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c02bff",
		x"f14000df40000070c160005fc160045fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2837fff",
		x"f080000840000071c0c0001140000072b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e05bff",
		x"f0a0001040000073c0e00041c0e00021b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e043ff",
		x"f100007f40000074c18001ffc18009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c241ffff",
		x"f0c0002040000075c1000041c10000c1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20083ff",
		x"f100008040000076b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200101",
		x"f0a0000fc1000057c10000d7c1000037c12000afc12001afc120006fc120016fc140003fc140023fc160017fc160057fc18001ffc18009ffc160037f",
		x"f0c0001fc10000b7c1000077c10000f7c12000efc12001efc120001fc120011fc140013fc140033fc160077fc16000ffc18005ffc1800dffc16004ff",
		x"f0c0003fc120009fc120019fc120005fc14000bfc14002bfc14001bfc14003bfc16002ffc16006ffc18003ffc1800bffc1a00fffc1a01fffc18007ff",
		x"f0a00007c0e00073c0e0000bc0e0004bc100009bc100005bc1200137c12000b7c140011fc140031fc160063fc160013fb0000000b0000000c160053f",
		x"f0c00017c10000dbc100003bc10000bbc12001b7c1200077c1200177c12000f7c140009fc160033fc180057fc1800d7fb0000000b0000000c160073f",
		x"f0c00037c100007bc10000fbc1000007c12001f7c120000fc120010fc140029fc16000bfc16004bfc180037fc1800b7fb0000000b0000000c16002bf",
		x"f0c0000fc1000087c1000047c10000c7c120008fc120018fc140019fc140039fc16006bfc16001bfc180077fc1800f7fb0000000b0000000c18000ff",
		x"f0e0005fc120004fc120014fc12000cfc140005fc140025fc140015fc16005bfc18008ffc18004ffc1a003ffc1a013ffb0000000b0000000c1800cff",
		x"f0e0003fc12001cfc120002fc120012fc140035fc14000dfc16003bfc16007bfc18002ffc1800affc1a00bffc1a01bffb0000000b0000000c1a007ff",
		x"f0c0002fc1000027c10000a7c1000067c12000afc12001afc14002dfc14001dfc160007fc160047fc18006ffc1800effb0000000b0000000c18001ff",
		x"f0e0007fc120006fc120016fc12000efc14003dfc140003fc160027fc160067fc18009ffc18005ffc1a017ffc1a00fffb0000000b0000000c1a01fff",
		x"f0a0000bc0e0007dc0e00003c0e00043c100003bc10000bbc12000cfc12001cfc16003bfc16007bfb0000000b0000000b0000000b0000000c160007f",
		x"f0a0001bc0e00023c0e00063c0e00013c100007bc10000fbc120002fc120012fc160047fc160027fb0000000b0000000b0000000b0000000c160067f",
		x"f0c0000fc0e00053c1000007c1000087c12000afc12001afc14000dfc14002dfc18002ffc1800affb0000000b0000000b0000000b0000000c18006ff",
		x"f0c0002fc1000047c10000c7c1000027c120006fc120016fc14001dfc14003dfc1800effc18001ffb0000000b0000000b0000000b0000000c18009ff",
		x"f0a00007c0c00015c0e00033c0e00073c10000a7c1000067c12000efc12001efc160017fc160057fb0000000b0000000b0000000b0000000c160037f",
		x"f0a00017c0e0000bc0e0004bc0e0002bc10000e7c1000017c120001fc120011fc160077fc16000ffb0000000b0000000b0000000b0000000c16004ff",
		x"f0c0001fc1000097c1000057c10000d7c120009fc120019fc140003fc140023fc18005ffc1800dffb0000000b0000000b0000000b0000000c18003ff",
		x"f0c0003fc1000037c10000b7c1000077c120005fc120015fc140013fc140033fc1800bffc18007ffb0000000b0000000b0000000b0000000c1800fff",
		x"f080000bc0a000194000007740000078c0e00043c0e00023c120018fc120004fb0000000b0000000b0000000b0000000b0000000b0000000c120014f",
		x"f0c00017c0c0003540000079c0e00063c100003bc10000bbc14002dfc14001dfb0000000b0000000b0000000b0000000b0000000b0000000c16001bf",
		x"f0c00037c0c0000d4000007ac0e00013c100007bc10000fbc14003dfc140003fb0000000b0000000b0000000b0000000b0000000b0000000c16005bf",
		x"f0e0004fc0e00053c1000007c1000087c12000cfc12001cfc16003bfc16007bfb0000000b0000000b0000000b0000000b0000000b0000000c1800aff",
		x"f0e0002fc0e00033c1000047c10000c7c120002fc120012fc160007fc160047fb0000000b0000000b0000000b0000000b0000000b0000000c18006ff",
		x"f0e0006fc0e00073c1000027c10000a7c12000afc12001afc160027fc160067fb0000000b0000000b0000000b0000000b0000000b0000000c1800eff",
		x"f0e0001fc0e0000bc1000067c10000e7c120006fc120016fc160017fc160057fb0000000b0000000b0000000b0000000b0000000b0000000c18001ff",
		x"f0800003c08000054000007bc0a0000dc0e00033c0e00073c12001efc140015fb0000000b0000000b0000000b0000000b0000000b0000000c140035f",
		x"f080000b4000007c4000007d4000007ec10000e7c1000017c14000dfc14002dfb0000000b0000000b0000000b0000000b0000000b0000000c160017f",
		x"f0a00007c0a0001d4000007f40000080c1000097c1000057c14001dfc160057fb0000000b0000000b0000000b0000000b0000000b0000000c160037f",
		x"f0c00017c0e0000bc10000d7c1000037c120001fc14003dfc180077fc1800f7fb0000000b0000000b0000000b0000000b0000000b0000000c1a005ff",
		x"f0e0001fc0e0004bc10000b7c1000077c140003fc140023fc18000ffc1a015ffb0000000b0000000b0000000b0000000b0000000b0000000c1a00dff",
		x"f0600005400000814000008240000083c100007bc12001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c140019f",
		x"f0a00003400000844000008540000086c140039fc140005fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16000bf",
		x"f0a000134000008740000088c0e0003bc140025fc140015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c180027f",
		x"f100003fc1200077c140035fc14000dfc1a00effc1a01effb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c00bff",
		x"f0600001400000894000008ac0800006c1000057c10000d7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c140003f",
		x"f0a0000bc080000e4000008bc0c0000dc140023fc140013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c180037f",
		x"f0c000074000008cc0e0001bc0e0005bc16003bfc1800b7fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a00dff",
		x"f0a0001bc08000014000008dc0c0002dc140033fc14000bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c180077f",
		x"f0a0000b4000008ec0c0002bc0c0001bc18004ffc1800cffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c013ff",
		x"f0a0001bc0800005c0c0003b4000008fc18002ffc1800affb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c033ff",
		x"f0a0000740000090c0c00007c0c00027c18006ffc1800effb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c00bff",
		x"f0e0001fc0c00017c100006f40000091c1c02bffc1c01bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2009fff",
		x"f060000640000092c080000cc0800002b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c140003f",
		x"f0c00017c080000ac0e0003bc0e0007bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a003ff",
		x"f0c00037c0800006c0e00007c0e00047b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18005ff",
		x"f120007fc0e00027c140023fc140013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e02fff",
		x"f0e0000fc080000ec0e00067c0e00017b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a013ff",
		x"f14001ffc0e00057c140033fc14000bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2007fff",
		x"f0600002400000934000009440000095b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16004ff",
		x"f0e0000740000096c1000017c12000f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e007ff",
		x"f06000024000009740000098c0a00009b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a003ff",
		x"f100008f40000099c120012fc14003afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2211fff",
		x"f100004f4000009ac12000afc140006fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2209fff",
		x"f08000044000009b4000009cc0c00011b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c01bff",
		x"f120001f4000009dc160025fc160065fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2607fff",
		x"f14002dfc0c00031c160015fc160055fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28b7fff",
		x"f14001dfc0c00009c160035fc160075fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2877fff",
		x"f08000044000009ec0c000314000009fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e03bff",
		x"f120003f400000a0c18000ffc1a009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c281ffff",
		x"f0a00008400000a1c0e00061c0e00011b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e023ff",
		x"f10000ffc0e00051c18005ffc1800dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c243ffff",
		x"f0c00010400000a2c1000021c10000a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20043ff",
		x"f1000040400000a3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200081",
		x"f0e0005fc0e0004bc1000017c1000097c12000efc12001efc160037fc160077fb0000000b0000000b0000000b0000000b0000000b0000000c18009ff",
		x"f0e0003fc0e0002bc1000057c10000d7c120001fc120011fc16000ffc16004ffb0000000b0000000b0000000b0000000b0000000b0000000c18005ff",
		x"f100007fc1000037c120009fc120019fc140023fc140013fc1800dffc18003ffb0000000b0000000b0000000b0000000b0000000b0000000c1a00fff",
		x"f10000ffc10000b7c120005fc120015fc140033fc14000bfc1800bffc18007ffb0000000b0000000b0000000b0000000b0000000b0000000c1a01fff",
		x"f0c00037c0c00003c0e0002bc0e0006bc120011fc120009fc18008ffc18004ffb0000000b0000000b0000000b0000000b0000000b0000000c1800cff",
		x"f0c0000fc0c00023c0e0001bc0e0005bc120019fc120005fc18002ffc1800affb0000000b0000000b0000000b0000000b0000000b0000000c18006ff",
		x"f0c0002fc0e0003bc10000f7c100000fc140013fc140033fc1800effc1a01dffb0000000b0000000b0000000b0000000b0000000b0000000c1a003ff",
		x"f0e0005fc0e0007bc100008fc100004fc14000bfc14002bfc18001ffc1a013ffb0000000b0000000b0000000b0000000b0000000b0000000c1a00bff",
		x"f0e0003fc0e00007c10000cfc100002fc14001bfc14003bfc18009ffc1a01bffb0000000b0000000b0000000b0000000b0000000b0000000c1a007ff",
		x"f0e0007fc0e00047c10000afc100006fc140007fc140027fc1a017ffc1a00fffb0000000b0000000b0000000b0000000b0000000b0000000c1a01fff",
		x"f0a0000bc0a0000b400000a4400000a5c1200177c14002dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16004bf",
		x"f0c0001b400000a6c10000fbc1000007c16002bfc16006bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a001ff",
		x"f0c0003b400000a7c1000087c1000047c16001bfc16005bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a011ff",
		x"f0c00007400000a8c10000c7c1000027c16003bfc16007bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a009ff",
		x"f0e00037c10000a7c12000f7c12001f7c1800a7fc180067fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c02bff",
		x"f0e00077c1000067c120000fc120010fc1800e7fc180017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c01bff",
		x"f0c00027400000a9c10000e7c1000017c160007fc160047fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a019ff",
		x"f0e0000fc1000097c120008fc120018fc180097fc180057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c03bff",
		x"f0800003c0600002400000aa400000abc120005fc120015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16007bf",
		x"f0c00027400000acc0c0001dc0c0003dc14002bfc160007fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a01dff",
		x"f0e0002fc0c00003c1000037c10000b7c1800f7fc18000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c017ff",
		x"f0e0006fc0c00023c1000077c10000f7c18008ffc18004ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c037ff",
		x"f0e0001f400000adc100000fc100008fc1800cffc18002ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c00fff",
		x"f0a00017c080000d400000ae400000afc18001ffc18009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c03bff",
		x"f100005fc0e00037c120009fc120019fc1e027ffc1e067ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2005fff",
		x"f0a0000fc0800003400000b0400000b1c18005ffc1800dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c007ff",
		x"f12001ffc120005fc160077fc16000ffc200dfffc221bfffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c243ffff",
		x"f0600001400000b2c0800001400000b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c14002bf",
		x"f0600006400000b4400000b5400000b6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16002ff",
		x"f0e00047400000b7c1000097c1000057b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e047ff",
		x"f0e00027400000b8c10000d7c12001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e027ff",
		x"f0e00067400000b9c1000037c120000fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e067ff",
		x"f0600006400000bac0a00019c0a00005b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a013ff",
		x"f10000cfc0a00015c140026fc140016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2219fff",
		x"f100002fc0a0000dc140036fc14000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2205fff",
		x"f10000afc0a0001dc14002efc14001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2215fff",
		x"f080000c400000bb400000bcc0c00029b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c03bff",
		x"f120011f400000bdc16000dfc16004dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2647fff",
		x"f120009f400000bec16002dfc16006dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2627fff",
		x"f080000c400000bfc0c00009400000c0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e07bff",
		x"f120013f400000c1c18008ffc1a019ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c289ffff",
		x"f12000bf400000c2c18004ffc1a005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c285ffff",
		x"f0a00018400000c3c0e00031c0e00071b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e063ff",
		x"f0c00030400000c4c1000061c10000e1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200c3ff",
		x"f10000c0400000c5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200181",
		x"f0e0004f400000c6c120004fc120014fc1800d7fc180037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c007ff",
		x"f0e0002fc1000057c12000cfc12001cfc1800b7fc180077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c027ff",
		x"f0e0006f400000c7c120002fc120012fc1800f7fc18000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c017ff",
		x"f0e0001fc10000d7c12000afc12001afc18008ffc18004ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c037ff",
		x"f0c00017400000c8c120006fc120016fc1800cffc18002ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c00fff",
		x"f0e0005fc1000037c12000efc12001efc1800affc18006ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c02fff",
		x"f0c00017400000c9c0e0003bc0e0007bc160047fc160027fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a003ff",
		x"f0c00037400000cac0e00007c0e00047c160067fc1800affb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a013ff",
		x"f0c0000fc0a00015c0e00027c0e00067c160017fc160057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a00bff",
		x"f10000ffc0e00017c12000dfc12001dfc1a01bffc1a007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e07fff",
		x"f10000dfc0e00077c120015fc12000dfc1e017ffc1e057ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2207fff",
		x"f100003fc0e0000fc12001dfc14003bfc1e037ffc1e077ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2217fff",
		x"f10000bfc0e0004fc120003fc120013fc1e00fffc1e04fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2003fff",
		x"f100007fc0e0002fc12000bfc140007fc1e02fffc1e06fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220ffff",
		x"f0800005400000cb400000cc400000cdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c14001bf",
		x"f0e0004f400000ce400000cfc1000077b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a00bff",
		x"f0800001400000d0400000d1c0a0000eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16006ff",
		x"f0e00017400000d2c10000b7c120010fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e017ff",
		x"f100004fc0a0001ec120008fc120018fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2002fff",
		x"f0e00057400000d3c1000077c120004fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e057ff",
		x"f10000cfc0a00001c120014fc12000cfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200afff",
		x"f100002fc0a00011c12001cfc120002fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e037ff",
		x"f0600001400000d4c0a00003400000d5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a00bff",
		x"f0800002400000d6400000d7c0c00019b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c007ff",
		x"f120019f400000d8c16001dfc16005dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2667fff",
		x"f120005f400000d9c16003dfc16007dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2617fff",
		x"f120015f400000dac160003fc160043fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2657fff",
		x"f0800002400000dbc0c00029c0e00015b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e007ff",
		x"f14001ffc0e00055c1800cffc1a015ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28dffff",
		x"f14003ffc0e00035c18002ffc1a00dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2afffff",
		x"f12001bfc0e00075c1800affc1a01dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2bfffff",
		x"f0a00004400000dcc0e00009c0e00049b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e013ff",
		x"f0c00008400000ddc1000011c1000091b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20023ff",
		x"f1000020400000deb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200041",
		x"f10000bfc120001fc14001dfc14003dfc1a005ffc1a015ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c01fff",
		x"f100007fc120011fc140003fc140023fc1a00dffc1a01dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e03fff",
		x"f10000ffc120009fc140013fc140033fc1a003ffc1a013ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e07fff",
		x"f0e0005fc0c00013c100004fc10000cfc18006ffc1800effb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c02fff",
		x"f0e0003fc0c00033c100002fc10000afc18001ffc18009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c01fff",
		x"f080000d400000dfc0a00009c0a00019b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c160037f",
		x"f0e0002fc0a00005c10000f7c100000fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a01bff",
		x"f100001fc0a00015c100008fc100004fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c007ff",
		x"f0e0006fc0a0000dc10000cfc100002fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c027ff",
		x"f14003ffc10000afc160077fc16000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200ffff",
		x"f0800009400000e0c0a00009c0a00019b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18001ff",
		x"f0e00037c0a00005c120012fc12000afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e077ff",
		x"f0e00077c0a00015c12001afc120006fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e00fff",
		x"f0e0000fc0a0000dc120016fc12000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e04fff",
		x"f0600005400000e1c0a00013400000e2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a01bff",
		x"f100006f400000e3c14003efc140001fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220dfff",
		x"f080000a400000e4400000e5c0c00039b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c027ff",
		x"f14003df400000e6c160023fc160063fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28f7fff",
		x"f140003f400000e7c160013fc160053fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c280ffff",
		x"f140023f400000e8c160033fc160073fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c288ffff",
		x"f140013f400000e9c16000bfc16004bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c284ffff",
		x"f0a0000a400000eac0c00019c0e0000db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e047ff",
		x"f0a00014400000ebc0e00029c0e00069b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e053ff",
		x"f0c00028400000ecc1000051c10000d1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200a3ff",
		x"f10000a0400000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200141",
		x"f0a00003400000eec0a0001d400000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16004ff",
		x"f0800005400000f0c0a0001d400000f1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18009ff",
		x"f0800003400000f2c0a0000b400000f3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a007ff",
		x"f12000ef400000f4c140021fc140011fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c241dfff",
		x"f12001ef400000f5c140031fc140009fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c243dfff",
		x"f0800006400000f6400000f7c0c00005b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c017ff",
		x"f140033f400000f8c16002bfc16006bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28cffff",
		x"f14000bfc0c00025c16001bfc16005bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c282ffff",
		x"f14002bfc0c00015c16003bfc16007bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28affff",
		x"f14001bfc0c00035c160007fc160047fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c286ffff",
		x"f14003bf400000f9c160027fc160067fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28effff",
		x"f0a0001a400000fac0c00039c0e0004db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e027ff",
		x"f0a0000c400000fbc0e00019c0e00059b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e033ff",
		x"f0c00018400000fcc1000031c10000b1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20063ff",
		x"f1000060400000fdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000c1",
		x"f0a00013400000fe400000ff40000100b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16002ff",
		x"f100009f40000101c12000efc12001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c017ff",
		x"f080000d40000102c0a0000340000103b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18005ff",
		x"f10000af40000104c12001efc140025fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2006fff",
		x"f080000b400001054000010640000107b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a017ff",
		x"f120001f40000108c140029fc160007fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2403fff",
		x"f120011f40000109c140019fc160047fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2423fff",
		x"f120009f4000010ac140039fc160027fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2413fff",
		x"f080000e4000010bc0c0000dc0c0002db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e037ff",
		x"f140007fc0c0001dc160017fc160057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c281ffff",
		x"f140027fc0c0003dc160037fc160077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c289ffff",
		x"f140017fc0c00003c16000ffc18004ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c285ffff",
		x"f0a000064000010cc0c00005c0e0002db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e067ff",
		x"f0a0001c4000010dc0e00039c0e00079b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e073ff",
		x"f0c000384000010ec1000071c10000f1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200e3ff",
		x"f10000e04000010fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001c1",
		x"f0a0000b40000110c0c00003c0c00023b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c16006ff",
		x"f100005f40000111c120001fc120011fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c037ff",
		x"f10000dfc0c00013c120009fc120019fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e06fff",
		x"f100003fc0c00033c120005fc120015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1c00fff",
		x"f0800003400001124000011340000114b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1800dff",
		x"f100006f40000115c120001fc140015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200efff",
		x"f10000ef40000116c120011fc140035fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2001fff",
		x"f0800007c02000004000011740000118b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1a00fff",
		x"f120019f40000119c140005fc140025fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2433fff",
		x"f120005f4000011ac140015fc160067fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c240bfff",
		x"f120015fc0c0001bc140035fc160017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c242bfff",
		x"f12000dfc0c0003bc14000dfc160057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c241bfff",
		x"f12001dfc0c00007c14002dfc160037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c243bfff",
		x"f08000014000011bc0c00023c0c00013b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e077ff",
		x"f0a000164000011cc0c00025c0e0006db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e017ff",
		x"f0a000024000011dc0e00005c0e00045b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e00bff",
		x"f0c000044000011ec1000009c1000089b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20013ff",
		x"f10000104000011fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200021",
		x"f0a0001bc0600000c0c0000b40000120b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1800dff",
		x"f10000bfc0c0002bc12000dfc12001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e01fff",
		x"f0a0000b4000012140000122c0c00013b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c18003ff",
		x"f100001f40000123c120009fc14000dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2009fff",
		x"f100009fc0c00033c14002dfc14001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2207fff",
		x"f100005fc0c0000bc14003dfc140003fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2005fff",
		x"f10000dfc0c0002bc140023fc140013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200dfff",
		x"f120003f40000124c14001dfc14003dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2407fff",
		x"f120013fc0c00027c140003fc160077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2427fff",
		x"f12000bf40000125c140023fc140013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2417fff",
		x"f12001bfc0c00017c140033fc16000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2437fff",
		x"f080000940000126c0c00033c0c0000bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e00fff",
		x"f0a0000e4000012740000128c0e0001db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e057ff",
		x"f0a0001240000129c0e00025c1000013b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e04bff",
		x"f0c000244000012ac1000049c10000c9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20093ff",
		x"f10000904000012bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200121",
		x"f120017f4000012cc14003bfc140007fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e05fff",
		x"f0a0001bc04000004000012dc0c0001bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1800bff",
		x"f100003f4000012ec140033fc14000bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2003fff",
		x"f10000bf4000012fc120019fc14002bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200bfff",
		x"f120007f40000130c14000bfc16004ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c240ffff",
		x"f120017f40000131c14002bfc16002ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c242ffff",
		x"f080000540000132c0c0002bc0c0001bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e04fff",
		x"f0a0001e4000013340000134c0e0005db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e037ff",
		x"f120007f40000135c18006ffc1a003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c283ffff",
		x"f0a0000a40000136c0e00065c1000093b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e02bff",
		x"f0c0001440000137c1000029c10000a9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20053ff",
		x"f100005040000138b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000a1",
		x"f12000ffc0e00037c140027fc140017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e03fff",
		x"f12000ffc0c0003bc14001bfc14003bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2217fff",
		x"f12001ffc0c00007c140007fc140027fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220ffff",
		x"f100007fc0c00027c140017fc140037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221ffff",
		x"f12000ffc0c00037c14001bfc16006ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c241ffff",
		x"f12001ffc0c0000fc14003bfc16001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c243ffff",
		x"f080000d40000139c0c0003b4000013ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e02fff",
		x"f0a000014000013bc0e0003dc0e0007db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e077ff",
		x"f120017fc0e00003c1800effc1a013ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28bffff",
		x"f12000ffc0e00043c18001ffc1a00bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c287ffff",
		x"f0a0001a4000013cc0e00015c1000053b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e06bff",
		x"f0c000344000013dc1000069c10000e9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200d3ff",
		x"f10000d04000013eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001a1",
		x"f08000034000013fc0c0000740000140b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e06fff",
		x"f140037f40000141c1800cffc18002ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28dffff",
		x"f0a0001140000142c0e00023c0e00063b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e00fff",
		x"f0a0000640000143c0e00055c10000d3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e01bff",
		x"f0c0000c40000144c1000019c1000099b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20033ff",
		x"f100003040000145b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200061",
		x"f080000b40000146c0c0002740000147b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e01fff",
		x"f14000ffc0e0000fc1800affc18006ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c283ffff",
		x"f14002ff40000148c1800effc18001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28bffff",
		x"f0a0000940000149c0e00013c0e00053b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2004fff",
		x"f0a000164000014ac0e00035c1000033b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e05bff",
		x"f0c0002c4000014bc1000059c10000d9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200b3ff",
		x"f10000b04000014cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200161",
		x"f08000074000014dc0c00017c0e0004fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e05fff",
		x"f14001ffc0e0002fc18009ffc18005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c287ffff",
		x"f14003ffc0e0006fc1800dffc18003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c28fffff",
		x"f0a000194000014ec0e00033c0e00073b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200cfff",
		x"f0a0000e4000014fc0e00075c10000b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e03bff",
		x"f0c0001c40000150c1000039c10000b9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20073ff",
		x"f100007040000151b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000e1",
		x"f0a0000fc0200000c0c00037c0e0001fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e03fff",
		x"f0a0000540000152c0e0000bc0e0004bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2002fff",
		x"f0a0001e40000153c0e0000dc1000073b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e07bff",
		x"f0c0003c40000154c1000079c10000f9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200f3ff",
		x"f10000f040000155b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001e1",
		x"f0a0001540000156c0e0002bc0e0006bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200afff",
		x"f0a0000140000157c0e0004dc10000f3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e007ff",
		x"f0c0000240000158c1000005c1000085b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2000bff",
		x"f100000840000159b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200011",
		x"f0a0000d4000015ac0e0001bc0e0005bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2006fff",
		x"f0a000114000015bc0e0002dc100000bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1e047ff",
		x"f0c000224000015cc1000045c10000c5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2008bff",
		x"f10000884000015db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200111",
		x"f0a0001d4000015ec0e0003bc0e0007bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200efff",
		x"f0c000094000015fc0e0006dc100008bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20027ff",
		x"f0c0001240000160c1000025c10000a5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2004bff",
		x"f100004840000161b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200091",
		x"f0a0000340000162c0e00007c0e00047b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2001fff",
		x"f0c0002940000163c0e0001dc100004bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200a7ff",
		x"f0c0003240000164c1000065c10000e5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200cbff",
		x"f10000c840000165b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200191",
		x"f0a0001340000166c0e00027c0e00067b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2009fff",
		x"f0c0001940000167c0e0005dc10000cbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20067ff",
		x"f0c0000a40000168c1000015c1000095b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2002bff",
		x"f100002840000169b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200051",
		x"f0a0000b4000016ac0e00017c0e00057b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2005fff",
		x"f0c000394000016bc0e0003dc100002bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200e7ff",
		x"f0c0002a4000016cc1000055c120006bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200abff",
		x"f10000a84000016db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200151",
		x"f0a0001b4000016ec0e00037c0e00077b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200dfff",
		x"f0c000054000016fc0e0007dc10000abb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20017ff",
		x"f0c0001a40000170c10000d5c120016bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2006bff",
		x"f100006840000171b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000d1",
		x"f0a0000740000172c0e0000fc0e0004fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2003fff",
		x"f0c0002540000173c0e00003c100006bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20097ff",
		x"f0c0003a40000174c1000035c12000ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200ebff",
		x"f10000e840000175b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001d1",
		x"f0a0001740000176c0e0002fc0e0006fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200bfff",
		x"f0c0001540000177c0e00043c10000ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20057ff",
		x"f0c0000640000178c10000b5c12001ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2001bff",
		x"f100001840000179b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200031",
		x"f0a0000f4000017ac0e0001fc0e0005fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2007fff",
		x"f0c000354000017bc0e00023c100001bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200d7ff",
		x"f0c000264000017cc1000075c120001bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2009bff",
		x"f10000984000017db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200131",
		x"f0c0001fc0200000c0e0003fc100007fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220ffff",
		x"f0c0000d4000017ec0e00063c100009bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20037ff",
		x"f0c000164000017fc10000f5c120011bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2005bff",
		x"f100005840000180b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000b1",
		x"f0c0002d40000181c100005bc10000dbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200b7ff",
		x"f0c0003640000182c100000dc120009bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200dbff",
		x"f10000d840000183b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001b1",
		x"f0c0001d40000184c100003bc10000bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20077ff",
		x"f0c0000e40000185c100008dc120019bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2003bff",
		x"f100003840000186b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200071",
		x"f0c0003d40000187c100007bc10000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200f7ff",
		x"f0c0002e40000188c100004dc120005bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200bbff",
		x"f10000b840000189b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200171",
		x"f0c000034000018ac1000007c1000087b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2000fff",
		x"f0c0001e4000018bc10000cdc120015bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2007bff",
		x"f10000784000018cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000f1",
		x"f0c000234000018dc1000047c10000c7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2008fff",
		x"f0c0003e4000018ec100002dc12000dbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200fbff",
		x"f10000f84000018fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001f1",
		x"f0c0001340000190c1000027c10000a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2004fff",
		x"f0c0000140000191c10000adc12001dbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20007ff",
		x"f100000440000192b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200009",
		x"f0c0003340000193c1000067c10000e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200cfff",
		x"f0c0002140000194c100006dc120003bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20087ff",
		x"f100008440000195b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200109",
		x"f0c0000b40000196c1000017c1000097b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2002fff",
		x"f0c0001140000197c10000edc120013bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20047ff",
		x"f100004440000198b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200089",
		x"f0c0002b40000199c1000057c10000d7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200afff",
		x"f0c000314000019ac100001dc12000bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200c7ff",
		x"f10000c44000019bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200189",
		x"f0c0001b4000019cc1000037c10000b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2006fff",
		x"f0c000094000019dc100009dc12001bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20027ff",
		x"f10000244000019eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200049",
		x"f0c0003b4000019fc1000077c10000f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200efff",
		x"f0c00029400001a0c100005dc120007bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200a7ff",
		x"f10000a4400001a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200149",
		x"f0c00007400001a2c100000fc100008fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2001fff",
		x"f0c00019400001a3c10000ddc120017bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20067ff",
		x"f1000064400001a4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000c9",
		x"f0c00027400001a5c100004fc10000cfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2009fff",
		x"f0c00039400001a6c100003dc12000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200e7ff",
		x"f10000e4400001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001c9",
		x"f0c00017400001a8c100002fc10000afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2005fff",
		x"f0c00005400001a9c10000bdc12001fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20017ff",
		x"f1000014400001aab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200029",
		x"f0c00037400001abc100006fc10000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200dfff",
		x"f0c00025400001acc100007dc1200007b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20097ff",
		x"f1000094400001adb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200129",
		x"f0c0000f400001aec100001fc100009fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2003fff",
		x"f0c00015400001afc10000fdc1200107b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c20057ff",
		x"f1000054400001b0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000a9",
		x"f0c0002f400001b1c100005fc10000dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c200bfff",
		x"f0e00035400001b2c1000003c1200087b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220d7ff",
		x"f10000d4400001b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001a9",
		x"f0c0001f400001b4c100003fc10000bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2007fff",
		x"f0e00075400001b5c1000083c1200187b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221d7ff",
		x"f1000034400001b6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200069",
		x"f0e0003fc0200000c100007fc12000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220ffff",
		x"f0e0000d400001b7c1000043c1200047b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c22037ff",
		x"f10000b4400001b8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200169",
		x"f0e0004d400001b9c10000c3c1200147b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c22137ff",
		x"f1000074400001bab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000e9",
		x"f0e0002d400001bbc1000023c12000c7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220b7ff",
		x"f10000f4400001bcb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001e9",
		x"f0e0006d400001bdc10000a3c12001c7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221b7ff",
		x"f100000c400001beb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200019",
		x"f0e0001d400001bfc1000063c1200027b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c22077ff",
		x"f100008c400001c0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200119",
		x"f0e0005d400001c1c10000e3c1200127b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c22177ff",
		x"f100004c400001c2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200099",
		x"f0e0003d400001c3c1000013c12000a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220f7ff",
		x"f10000cc400001c4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200199",
		x"f0e0007d400001c5c1000093c12001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221f7ff",
		x"f100002c400001c6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200059",
		x"f0e00003400001c7c1000053c1200067b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2200fff",
		x"f10000ac400001c8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200159",
		x"f0e00043400001c9c10000d3c1200167b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2210fff",
		x"f100006c400001cab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000d9",
		x"f0e00023400001cbc1000033c12000e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2208fff",
		x"f10000ec400001ccb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001d9",
		x"f0e00063400001cdc10000b3c12001e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2218fff",
		x"f100001c400001ceb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200039",
		x"f0e00013400001cfc1000073c1200017b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2204fff",
		x"f100009c400001d0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200139",
		x"f0e00053400001d1c10000f3c1200117b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2214fff",
		x"f100005c400001d2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000b9",
		x"f0e00033400001d3c100000bc1200097b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220cfff",
		x"f10000dc400001d4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001b9",
		x"f0e00073400001d5c100008bc1200197b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221cfff",
		x"f100003c400001d6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200079",
		x"f0e0000b400001d7c100004bc1200057b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2202fff",
		x"f10000bc400001d8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200179",
		x"f0e0004b400001d9c10000cbc1200157b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2212fff",
		x"f100007c400001dab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000f9",
		x"f0e0002b400001dbc100002bc12000d7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220afff",
		x"f10000fc400001dcb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001f9",
		x"f0e0006b400001ddc10000abc12001d7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221afff",
		x"f1000002400001deb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200005",
		x"f0e0001b400001dfc1200037c1200137b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2206fff",
		x"f1000082400001e0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200105",
		x"f0e0005b400001e1c12000b7c12001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2216fff",
		x"f1000042400001e2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200085",
		x"f0e0003b400001e3c1200077c1200177b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220efff",
		x"f10000c2400001e4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200185",
		x"f0e0007b400001e5c12000f7c12001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221efff",
		x"f1000022400001e6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200045",
		x"f0e00007400001e7c120000fc120010fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2201fff",
		x"f10000a2400001e8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200145",
		x"f0e00047400001e9c120008fc120018fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2211fff",
		x"f1000062400001eab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000c5",
		x"f0e00027400001ebc120004fc120014fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2209fff",
		x"f10000e2400001ecb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001c5",
		x"f0e00067400001edc12000cfc12001cfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2219fff",
		x"f1000012400001eeb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200025",
		x"f0e00017400001efc120002fc120012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2205fff",
		x"f1000092400001f0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200125",
		x"f0e00057400001f1c12000afc12001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2215fff",
		x"f1000052400001f2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000a5",
		x"f0e00037400001f3c120006fc120016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220dfff",
		x"f10000d2400001f4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001a5",
		x"f0e00077400001f5c12000efc12001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221dfff",
		x"f1000032400001f6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200065",
		x"f0e0000f400001f7c120001fc120011fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2203fff",
		x"f10000b2400001f8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200165",
		x"f0e0004f400001f9c120009fc120019fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2213fff",
		x"f1000072400001fab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000e5",
		x"f0e0002f400001fbc120005fc120015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220bfff",
		x"f10000f2400001fcb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001e5",
		x"f0e0006f400001fdc12000dfc12001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221bfff",
		x"f100000a400001feb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200015",
		x"f0e0001f400001ffc120003fc120013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2207fff",
		x"f100008a40000200b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200115",
		x"f0e0005f40000201c12000bfc12001bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c2217fff",
		x"f100004a40000202b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200095",
		x"f0e0003f40000203c120007fc120017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c220ffff",
		x"f10000ca40000204b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200195",
		x"f0e0007fc0200000c12000ffc14001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c221ffff",
		x"f100002a40000205b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200055",
		x"f10000aa40000206b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200155",
		x"f100006a40000207b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000d5",
		x"f10000ea40000208b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001d5",
		x"f100001a40000209b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200035",
		x"f100009a4000020ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200135",
		x"f100005a4000020bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000b5",
		x"f10000da4000020cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001b5",
		x"f100003a4000020db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200075",
		x"f10000ba4000020eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200175",
		x"f100007a4000020fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000f5",
		x"f10000fa40000210b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001f5",
		x"f100000640000211b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120000d",
		x"f100008640000212b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120010d",
		x"f100004640000213b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120008d",
		x"f10000c640000214b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120018d",
		x"f100002640000215b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120004d",
		x"f10000a640000216b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120014d",
		x"f100006640000217b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000cd",
		x"f10000e640000218b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001cd",
		x"f100001640000219b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120002d",
		x"f10000964000021ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120012d",
		x"f10000564000021bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000ad",
		x"f10000d64000021cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001ad",
		x"f10000364000021db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120006d",
		x"f10000b64000021eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120016d",
		x"f10000764000021fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000ed",
		x"f10000f640000220b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001ed",
		x"f100000e40000221b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120001d",
		x"f100008e40000222b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120011d",
		x"f100004e40000223b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120009d",
		x"f10000ce40000224b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120019d",
		x"f100002e40000225b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120005d",
		x"f10000ae40000226b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120015d",
		x"f100006e40000227b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000dd",
		x"f10000ee40000228b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001dd",
		x"f100001e40000229b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120003d",
		x"f100009e4000022ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120013d",
		x"f100005e4000022bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000bd",
		x"f10000de4000022cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001bd",
		x"f100003e4000022db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120007d",
		x"f10000be4000022eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120017d",
		x"f100007e4000022fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000fd",
		x"f10000fe40000230b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001fd",
		x"f100000140000231b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200003",
		x"f100008140000232b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200103",
		x"f100004140000233b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200083",
		x"f10000c140000234b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200183",
		x"f100002140000235b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200043",
		x"f10000a140000236b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200143",
		x"f100006140000237b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000c3",
		x"f10000e140000238b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001c3",
		x"f100001140000239b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200023",
		x"f10000914000023ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200123",
		x"f10000514000023bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000a3",
		x"f10000d14000023cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001a3",
		x"f10000314000023db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200063",
		x"f10000b14000023eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200163",
		x"f10000714000023fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000e3",
		x"f10000f140000240b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001e3",
		x"f100000940000241b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200013",
		x"f100008940000242b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200113",
		x"f100004940000243b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200093",
		x"f10000c940000244b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200193",
		x"f100002940000245b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200053",
		x"f10000a940000246b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200153",
		x"f100006940000247b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000d3",
		x"f10000e940000248b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001d3",
		x"f100001940000249b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200033",
		x"f10000994000024ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200133",
		x"f10000594000024bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000b3",
		x"f10000d94000024cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001b3",
		x"f10000394000024db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200073",
		x"f10000b94000024eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200173",
		x"f10000794000024fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000f3",
		x"f10000f940000250b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001f3",
		x"f100000540000251b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120000b",
		x"f100008540000252b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120010b",
		x"f100004540000253b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120008b",
		x"f10000c540000254b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120018b",
		x"f100002540000255b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120004b",
		x"f10000a540000256b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120014b",
		x"f100006540000257b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000cb",
		x"f10000e540000258b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001cb",
		x"f100001540000259b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120002b",
		x"f10000954000025ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120012b",
		x"f10000554000025bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000ab",
		x"f10000d54000025cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001ab",
		x"f10000354000025db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120006b",
		x"f10000b54000025eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120016b",
		x"f10000754000025fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000eb",
		x"f10000f540000260b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001eb",
		x"f100000d40000261b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120001b",
		x"f100008d40000262b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120011b",
		x"f100004d40000263b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120009b",
		x"f10000cd40000264b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120019b",
		x"f100002d40000265b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120005b",
		x"f10000ad40000266b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120015b",
		x"f100006d40000267b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000db",
		x"f10000ed40000268b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001db",
		x"f100001d40000269b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120003b",
		x"f100009d4000026ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120013b",
		x"f100005d4000026bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000bb",
		x"f10000dd4000026cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001bb",
		x"f100003d4000026db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120007b",
		x"f10000bd4000026eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120017b",
		x"f100007d4000026fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000fb",
		x"f10000fd40000270b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001fb",
		x"f100000340000271b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200007",
		x"f100008340000272b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200107",
		x"f100004340000273b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200087",
		x"f10000c340000274b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200187",
		x"f100002340000275b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200047",
		x"f10000a340000276b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200147",
		x"f100006340000277b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000c7",
		x"f10000e340000278b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001c7",
		x"f100001340000279b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200027",
		x"f10000934000027ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200127",
		x"f10000534000027bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000a7",
		x"f10000d34000027cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001a7",
		x"f10000334000027db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200067",
		x"f10000b34000027eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200167",
		x"f10000734000027fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000e7",
		x"f10000f340000280b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001e7",
		x"f100000b40000281b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200017",
		x"f100008b40000282b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200117",
		x"f100004b40000283b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200097",
		x"f10000cb40000284b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200197",
		x"f100002b40000285b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200057",
		x"f10000ab40000286b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200157",
		x"f100006b40000287b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000d7",
		x"f10000eb40000288b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001d7",
		x"f100001b40000289b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200037",
		x"f100009b4000028ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200137",
		x"f100005b4000028bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000b7",
		x"f10000db4000028cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001b7",
		x"f100003b4000028db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200077",
		x"f10000bb4000028eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c1200177",
		x"f100007b4000028fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000f7",
		x"f10000fb40000290b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001f7",
		x"f100000740000291b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120000f",
		x"f100008740000292b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120010f",
		x"f100004740000293b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120008f",
		x"f10000c740000294b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120018f",
		x"f100002740000295b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120004f",
		x"f10000a740000296b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120014f",
		x"f100006740000297b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000cf",
		x"f10000e740000298b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001cf",
		x"f100001740000299b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120002f",
		x"f10000974000029ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120012f",
		x"f10000574000029bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000af",
		x"f10000d74000029cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001af",
		x"f10000374000029db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120006f",
		x"f10000b74000029eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120016f",
		x"f10000774000029fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000ef",
		x"f10000f7400002a0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001ef",
		x"f100000f400002a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120001f",
		x"f100008f400002a2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120011f",
		x"f100004f400002a3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120009f",
		x"f10000cf400002a4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120019f",
		x"f100002f400002a5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120005f",
		x"f10000af400002a6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120015f",
		x"f100006f400002a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000df",
		x"f10000ef400002a8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001df",
		x"f100001f400002a9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120003f",
		x"f100009f400002aab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120013f",
		x"f100005f400002abb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000bf",
		x"f10000df400002acb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001bf",
		x"f100003f400002adb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120007f",
		x"f10000bf400002aeb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c120017f",
		x"f100007f400002afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12000ff",
		x"f10000ffc0200000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c12001ff"
    );
end ccsds_constants;

package body ccsds_constants is
	
end ccsds_constants;
