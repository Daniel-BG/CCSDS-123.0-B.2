----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02.03.2021 10:35:20
-- Design Name: 
-- Module Name: constants - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.ccsds_math_functions.all;

package ccsds_constants is
	--IMAGE CONSTANTS
	type local_sum_t is (WIDE_NEIGHBOR_ORIENTED, WIDE_COLUMN_ORIENTED);
	type relocation_mode_t is (VERTICAL_TO_DIAGONAL, DIAGONAL_TO_VERTICAL); 
	
	--OTHER CONSTANTS
	constant STDLV_ONE: std_logic_vector(0 downto 0) := "1";
	constant STDLV_ZERO: std_logic_vector(0 downto 0) := "0";
	
	--FIXED CONSTANTS
	constant CONST_TINC_MIN				: integer := 4;
	constant CONST_TINC_MAX				: integer := 11;
	constant CONST_TINC_BITS 			: integer := 4;
	constant CONST_VMIN					: integer := -6;
	constant CONST_VMAX					: integer := 9;
	constant CONST_VMINMAX_BITS 		: integer := 5;
	constant CONST_WEO_MIN				: integer := -6;
	constant CONST_WEO_MAX				: integer := 5;
	constant CONST_WEO_BITS 			: integer := 4;
	constant CONST_MAX_RES_VAL 			: integer := 4;
	constant CONST_DATA_WIDTH_MAX		: integer := 32;
	constant CONST_DATA_WIDTH_MIN		: integer := 2;
	constant CONST_OMEGA_WIDTH_MAX		: integer := 19;
	constant CONST_OMEGA_WIDTH_MIN		: integer := 4;
	constant CONST_WUSE_BITS 			: integer := 7;

	--CONSTANTS THAT CAN ALTER RESOURCE USE
	constant CONST_MAX_DATA_WIDTH		: integer := 16;				--maximum allowed bits for inputs (Can be set lower through cfg ports)
	constant CONST_MAX_OMEGA			: integer := 19;				--maximum allowed bits for weights (Can be set lower through cfg ports)
	constant CONST_MIN_OMEGA			: integer := 4;
	constant CONST_MAX_P				: integer := 3;					--maximum allowed bits for previous bands used in prediction
	constant CONST_MAX_BANDS			: integer := 256;				--maximum allowed size in the x direction (Can be set lower through cfg ports)
	constant CONST_MAX_LINES			: integer := 1024;				--maximum allowed size in the y direction (Can be set lower through cfg ports)
	constant CONST_MAX_SAMPLES			: integer := 512;  				--maximum allowed size in the z direction (Can be set lower through cfg ports)
	
	--DERIVED CONSTANTS
	constant CONST_MAX_SAMPLES_PER_BAND	: integer := CONST_MAX_SAMPLES * CONST_MAX_LINES;
	
	constant CONST_MAX_X_VALUE			: integer := CONST_MAX_SAMPLES - 1;	--maximum allowed size in the x direction (Can be set lower through cfg ports)
	constant CONST_MAX_Y_VALUE			: integer := CONST_MAX_LINES - 1;	--maximum allowed size in the y direction (Can be set lower through cfg ports)
	constant CONST_MAX_Z_VALUE			: integer := CONST_MAX_BANDS - 1;  	--maximum allowed size in the z direction (Can be set lower through cfg ports)
	constant CONST_MAX_T_VALUE			: integer := CONST_MAX_SAMPLES_PER_BAND - 1;
	
	constant CONST_ABS_ERR_BITS 		: integer := MIN(CONST_MAX_DATA_WIDTH - 1, 16); 
	constant CONST_REL_ERR_BITS 		: integer := MIN(CONST_MAX_DATA_WIDTH - 1, 16); 
	
	constant CONST_MAX_WEIGHT_BITS		: integer := CONST_MAX_OMEGA + 3;
	constant CONST_MAX_C				: integer := CONST_MAX_P + 3; --number of previous bands plus 3 (full pred mode)
	constant CONST_MAX_OMEGA_WIDTH_BITS	: integer := BITS(CONST_MAX_OMEGA);		
	constant CONST_MAX_DATA_WIDTH_BITS	: integer := BITS(CONST_MAX_DATA_WIDTH);	
	constant CONST_MAX_P_WIDTH_BITS  	: integer := BITS(CONST_MAX_P);
	constant CONST_MAX_C_BITS			: integer := BITS(CONST_MAX_C);
	
	constant CONST_MAX_X_VALUE_BITS		: integer := BITS(CONST_MAX_X_VALUE);
	constant CONST_MAX_Y_VALUE_BITS		: integer := BITS(CONST_MAX_Y_VALUE);
	constant CONST_MAX_Z_VALUE_BITS		: integer := BITS(CONST_MAX_Z_VALUE);
	constant CONST_MAX_T_VALUE_BITS		: integer := BITS(CONST_MAX_T_VALUE);
	
	constant CONST_MAX_BANDS_BITS		: integer := BITS(CONST_MAX_BANDS);
	constant CONST_MAX_LINES_BITS		: integer := BITS(CONST_MAX_LINES);
	constant CONST_MAX_SAMPLES_BITS		: integer := BITS(CONST_MAX_SAMPLES);
	
	constant CONST_CQBC_BITS			: integer := CONST_MAX_DATA_WIDTH;
	constant CONST_QI_BITS				: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_LSUM_BITS			: integer := CONST_MAX_DATA_WIDTH + 2;
	constant CONST_LDIF_BITS			: integer := CONST_MAX_DATA_WIDTH + 3;
	constant CONST_DRSR_BITS 			: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_DRPSV_BITS 			: integer := CONST_MAX_DATA_WIDTH + 1;
	constant CONST_DRPE_BITS 			: integer := CONST_MAX_DATA_WIDTH + 2;
	constant CONST_PR_BITS 				: integer := CONST_MAX_DATA_WIDTH + 1;
	
	constant CONST_MEV_BITS 			: integer := MAX(CONST_ABS_ERR_BITS, CONST_REL_ERR_BITS);
	constant CONST_PCLD_BITS 			: integer := CONST_MAX_WEIGHT_BITS + BITS((2**CONST_MAX_DATA_WIDTH - 1)*(8*CONST_MAX_P + 19));
	constant CONST_HRPSV_BITS			: integer := CONST_MAX_OMEGA + 2 + CONST_MAX_DATA_WIDTH; 
	
	constant CONST_RES_BITS				: integer := BITS(CONST_MAX_RES_VAL);
	constant CONST_DAMPING_BITS			: integer := CONST_MAX_RES_VAL;
	constant CONST_OFFSET_BITS			: integer := CONST_MAX_RES_VAL;
	
	constant CONST_DIFFVEC_BITS 		: integer := CONST_MAX_C * CONST_LDIF_BITS;
	constant CONST_CLDVEC_BITS 			: integer := CONST_MAX_P * CONST_LDIF_BITS;
	constant CONST_DIRDIFFVEC_BITS		: integer := 3 * CONST_LDIF_BITS;
	constant CONST_WEIGHTVEC_BITS		: integer := CONST_MAX_C * CONST_MAX_WEIGHT_BITS;
	
	constant CONST_W_UPDATE_BITS		: integer := CONST_LDIF_BITS - CONST_VMIN - CONST_WEO_MIN - CONST_DATA_WIDTH_MIN + CONST_OMEGA_WIDTH_MAX; --should be 64
	
	constant CONST_THETA_BITS			: integer := CONST_MAX_DATA_WIDTH;
	constant CONST_MQI_BITS				: integer := CONST_MAX_DATA_WIDTH;
	
	--ENCODER CONSTANTS
	constant CONST_MIN_GAMMA_ZERO		: integer := 1;
	constant CONST_MAX_GAMMA_ZERO		: integer := 8;
	constant CONST_MAX_GAMMA_STAR		: integer := 11;
	constant CONST_MAX_COUNTER_BITS 	: integer := CONST_MAX_GAMMA_STAR;
	constant CONST_MAX_ACC_BITS			: integer := CONST_MAX_GAMMA_STAR + CONST_MAX_DATA_WIDTH;
	constant CONST_MAX_HR_ACC_BITS		: integer := CONST_MAX_ACC_BITS + 2;
	constant CONST_MAX_K				: integer := CONST_MAX_DATA_WIDTH - 2;
	constant CONST_MAX_K_BITS			: integer := BITS(CONST_MAX_K);
	constant CONST_U_MAX_MIN			: integer := 8;
	constant CONST_U_MAX_MAX			: integer := 32;
	constant CONST_U_MAX_BITS			: integer := BITS(CONST_U_MAX_MAX);
	
	constant CONST_MAX_CODE_LENGTH		: integer := CONST_U_MAX_MAX + CONST_MAX_DATA_WIDTH;
	constant CONST_MAX_CODE_LENGTH_BITS : integer := BITS(CONST_MAX_CODE_LENGTH);
	
	constant CONST_OUTPUT_CODE_LENGTH 	: integer := 64;
	constant CONST_OUTPUT_CODE_LENGTH_BITS: integer := 7;
	
	
	subtype threshold_value_t is std_logic_vector (18 downto 0);
    type threshold_table_t is array (0 to 15) of threshold_value_t;

    constant CONST_THRESHOLD_TABLE : threshold_table_t := (
		x"4A0E8",
		x"3707C",
		x"28C43",
		x"1F6A0",
		x"1756D",
		x"11026",
		x"0C5F6",
		x"08852",
		x"05B23",
		x"03A57",
		x"02442",
		x"01586",
		x"00C7B",
		x"00788",
		x"00458",
		x"00198"
	);
	
	type input_symbol_limit_t is array (0 to 15) of std_logic_vector(3 downto 0);
	constant CONST_INPUT_SYMBOL_LIMIT : input_symbol_limit_t := (
		x"C", x"A", x"8", x"6",
		x"6", x"4", x"4", x"4",
		x"2", x"2", x"2", x"2",
		x"0", x"0", x"0", x"0"		
	);
	
	constant CONST_INPUT_SYMBOL_X: std_logic_vector := "1101";
	
	constant CONST_CODEWORD_BITS: integer := 21;
	constant CONST_CODEWORD_LENGTH_BITS: integer := 5;
	
	constant CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT: integer := 688;
	constant CONST_LOW_ENTROPY_CODING_TABLE_ADDRESS_BITS: integer := bits(CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT);
	
	subtype bin_table_t is std_logic_vector (32*15-1 downto 0);
    type table_rom_t is array (0 to CONST_LOW_ENTROPY_CODING_TABLE_AMOUNT - 1) of bin_table_t;

    constant CONST_LOW_ENTROPY_CODING_TABLE : table_rom_t := (
		x"f000002040000010c0000060c0000064c000006240000011c0000086c000008e4000001240000013c00000a1c00000b1c00000c5c00000e5c00000a9",
		x"f0000020400000144000001540000016c0000060c0000064c0000082c000008ac00000a6c00000b6c00000cd40000017b0000000b0000000c00000ed",
		x"f0000020c00000404000001840000019c0000062c00000664000001a4000001bc00000d9c00000f9b0000000b0000000b0000000b0000000c00000c5",
		x"f00000204000001cc00000404000001d4000001e4000001fc00000ae40000020b0000000b0000000b0000000b0000000b0000000b0000000c00000c5",
		x"f000002040000021c0000040c0000042c0000081c0000089c00000f3c00000f3b0000000b0000000b0000000b0000000b0000000b0000000c0000127",
		x"f0000020c0000020c000004140000022c00000a3c00000b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00000fb",
		x"f000004040000023400000244000002540000026c00000ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00000204000002740000028c000006140000029c00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000404000002a4000002b4000002cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00000604000002dc0000082c000008ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000015f",
		x"f00000604000002e4000002fc00000a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f000008040000030c00000a140000031b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f000008040000032c00000c1c00000e1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f00000a04000003340000034c00000e1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000c040000035c0000101c0000181b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f000010040000036b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000121",
		x"f0000041c00000b94000003740000038c00000d5c00000f5c00000cdc00000edc00000f3c00000f3c000013bc00001bbc000012fc000012fc000017b",
		x"f0000063c00000ddc00000fdc00000c3c00000e340000039c00000f3c00000f3c00001fbc0000107c00001afc00001afc000016fc000016fc0000187",
		x"f00000a7c00000ebc00000ebc00000ebc0000147c00001c7c0000127c00001a7c00001efc00001efc000015fc000035fc000017fc000057fc00001df",
		x"f00000b7c00000ebc00000fbc00000fbc0000167c00001e7c0000117c0000197c000012fc000012fc00003dfc00001dfc000037fc000077fc00003df",
		x"f00000614000003ac00000aec00000be4000003b4000003cc00000ddc00000fdc00000f3c00000f3c00001e7c00001e7b0000000b0000000c000012b",
		x"f0000065c00000a1c00000b1c00000a94000003dc00000c34000003e4000003fc00001abc000016bc0000137c0000137b0000000b0000000c00001b7",
		x"f0000063c00000b9c00000a5c00000b540000040c00000e340000041c00000f3c00001ebc000011bc00001b7c0000177b0000000b0000000c0000177",
		x"f00000ffc00001f7c00001f7c0000137c00001efc00003efc000015fc000035fc000037fc00001ffc0000dffc0001dffb0000000b0000000c00009ff",
		x"f0000061c000008140000042400000434000004440000045c00000f5c00000f5c000016bc00001f7b0000000b0000000b0000000b0000000c00001f7",
		x"f00000654000004640000047c00000a94000004840000049c00000edc00000edc00001ebc000012fb0000000b0000000b0000000b0000000c000012f",
		x"f00000a3c00000e5c00000edc00000edc000011bc000019bc00001afc00001afc00001ffc00005ffb0000000b0000000b0000000b0000000c00003ff",
		x"f00000b3c00000fdc00000fdc00000fdc000015bc00001dbc000016fc000016fc00007ffc00001ffb0000000b0000000b0000000b0000000c00005ff",
		x"f00000614000004ac0000082c000008ac00000bec00000a1c00000edc00000edb0000000b0000000b0000000b0000000b0000000b0000000c000016b",
		x"f0000065c00000864000004b4000004c4000004dc00000e5c00001ebc000011bb0000000b0000000b0000000b0000000b0000000b0000000c000019b",
		x"f0000083c00000b14000004e4000004fc00000fdc00000fdc0000177c0000177b0000000b0000000b0000000b0000000b0000000b0000000c00001f7",
		x"f00000a7c00000a940000050c00000d5c00000fdc00000fdc00001f7c000012fb0000000b0000000b0000000b0000000b0000000b0000000c00001df",
		x"f00000efc00000e3c000015bc00001dbc000012fc00001afc00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000414000005140000052400000534000005440000055c00001a7c0000167b0000000b0000000b0000000b0000000b0000000b0000000c00001ef",
		x"f0000061400000564000005740000058c00000fb40000059b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b7",
		x"f00000424000005ac00000604000005bc00000ebc00000ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f0000085c00000644000005cc00000a9c00001efc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f000008d4000005dc00000b9c00000a5c000013fc000013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f000017fc00000ebc00001bfc00001bfc00005ffc00015ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f0000041c00000204000005e4000005fc00001efc000013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000037f",
		x"f00000834000006040000061c00000cbc000077fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00001ffc000013fc000057fc000037fc0001fffc000bfffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f00000624000006240000063c0000084b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00000c74000006440000065c00000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000e74000006640000067c00000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00009ff",
		x"f000006440000068c000008640000069b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000644000006a4000006bc00000b1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000dff",
		x"f000010f4000006cc000012fc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00000884000006d4000006e4000006fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002bff",
		x"f00001df40000070c000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0037fff",
		x"f000008840000071c00000d140000072b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005bff",
		x"f00000b040000073c00000e1c00000e1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00043ff",
		x"f000017f40000074c00001ffc00009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f00000e040000075c0000141c00001c1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00083ff",
		x"f000018040000076b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000121",
		x"f00000afc0000157c00001d7c0000137c00001afc00001afc000016fc000016fc000017fc000037fc000017fc000057fc00001ffc00009ffc000037f",
		x"f00000dfc00001b7c0000177c00001f7c00001efc00001efc000013fc000013fc000017fc000037fc000077fc00001ffc00005ffc0000dffc00005ff",
		x"f00000ffc00001bfc00001bfc000017fc00001ffc00003ffc00001ffc00003ffc00003ffc00007ffc00003ffc0000bffc0000fffc0001fffc00007ff",
		x"f00000a7c00000f3c00000ebc00000ebc000019bc000015bc0000137c00001b7c000015fc000035fc000077fc000017fb0000000b0000000c000057f",
		x"f00000d7c00001dbc000013bc00001bbc00001b7c0000177c0000177c00001f7c00001dfc000037fc00005ffc0000dffb0000000b0000000c000077f",
		x"f00000f7c000017bc00001fbc0000107c00001f7c000012fc000012fc00003dfc00001ffc00005ffc00003ffc0000bffb0000000b0000000c00003ff",
		x"f00000cfc0000187c0000147c00001c7c00001afc00001afc00001dfc00003dfc00007ffc00001ffc00007ffc0000fffb0000000b0000000c00001ff",
		x"f00000ffc000016fc000016fc00001efc000015fc000035fc000015fc00005ffc00009ffc00005ffc00003ffc00013ffb0000000b0000000c0000dff",
		x"f00000ffc00001efc000012fc000012fc000035fc00001dfc00003ffc00007ffc00003ffc0000bffc0000bffc0001bffb0000000b0000000c00007ff",
		x"f00000efc0000127c00001a7c0000167c00001afc00001afc00003dfc00001dfc000017fc000057fc00007ffc0000fffb0000000b0000000c00001ff",
		x"f00000ffc000016fc000016fc00001efc00003dfc000017fc000037fc000077fc00009ffc00005ffc00017ffc0000fffb0000000b0000000c0001fff",
		x"f00000abc00000fdc00000e3c00000e3c000013bc00001bbc00001efc00001efc00003ffc00007ffb0000000b0000000b0000000b0000000c000017f",
		x"f00000bbc00000e3c00000e3c00000f3c000017bc00001fbc000012fc000012fc000057fc000037fb0000000b0000000b0000000b0000000c000077f",
		x"f00000cfc00000f3c0000107c0000187c00001afc00001afc00001dfc00003dfc00003ffc0000bffb0000000b0000000b0000000b0000000c00007ff",
		x"f00000efc0000147c00001c7c0000127c000016fc000016fc00001dfc00003dfc0000fffc00001ffb0000000b0000000b0000000b0000000c00009ff",
		x"f00000a7c00000d5c00000f3c00000f3c00001a7c0000167c00001efc00001efc000017fc000057fb0000000b0000000b0000000b0000000c000037f",
		x"f00000b7c00000ebc00000ebc00000ebc00001e7c0000117c000013fc000013fc000077fc00001ffb0000000b0000000b0000000b0000000c00005ff",
		x"f00000dfc0000197c0000157c00001d7c00001bfc00001bfc000017fc000037fc00005ffc0000dffb0000000b0000000b0000000b0000000c00003ff",
		x"f00000ffc0000137c00001b7c0000177c000017fc000017fc000017fc000037fc0000bffc00007ffb0000000b0000000b0000000b0000000c0000fff",
		x"f000008bc00000b94000007740000078c00000e3c00000e3c00001afc000016fb0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00000d7c00000f540000079c00000e3c000013bc00001bbc00003dfc00001dfb0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000f7c00000cd4000007ac00000f3c000017bc00001fbc00003dfc000017fb0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f00000efc00000f3c0000107c0000187c00001efc00001efc00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f00000efc00000f3c0000147c00001c7c000012fc000012fc000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000efc00000f3c0000127c00001a7c00001afc00001afc000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000ffc00000ebc0000167c00001e7c000016fc000016fc000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f0000083c00000854000007bc00000adc00000f3c00000f3c00001efc000015fb0000000b0000000b0000000b0000000b0000000b0000000c000035f",
		x"f000008b4000007c4000007d4000007ec00001e7c0000117c00001dfc00003dfb0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f00000a7c00000bd4000007f40000080c0000197c0000157c00001dfc000057fb0000000b0000000b0000000b0000000b0000000b0000000c000037f",
		x"f00000d7c00000ebc00001d7c0000137c000013fc00003dfc00007ffc0000fffb0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f00000ffc00000ebc00001b7c0000177c000017fc000037fc00001ffc00015ffb0000000b0000000b0000000b0000000b0000000b0000000c0000dff",
		x"f0000065400000814000008240000083c000017bc00001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001df",
		x"f00000a3400000844000008540000086c00003dfc000015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000b34000008740000088c00000fbc000035fc000015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f000013fc0000177c000035fc00001dfc0000fffc0001fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f0000061400000894000008ac0000086c0000157c00001d7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f00000abc000008e4000008bc00000cdc000037fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000c74000008cc00000fbc00000fbc00003ffc0000bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000dff",
		x"f00000bbc00000814000008dc00000edc000037fc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000ab4000008ec00000ebc00000dbc00005ffc0000dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00013ff",
		x"f00000bbc0000085c00000fb4000008fc00003ffc0000bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00033ff",
		x"f00000a740000090c00000c7c00000e7c00007ffc0000fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f00000ffc00000d7c000016f40000091c0002bffc0001bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009fff",
		x"f000006640000092c000008cc0000082b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f00000d7c000008ac00000fbc00000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000f7c0000086c00000e7c00000e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f000017fc00000e7c000037fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000efc000008ec00000e7c00000f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00013ff",
		x"f00001ffc00000f7c000037fc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f0000062400000934000009440000095b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f00000e740000096c0000117c00001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000624000009740000098c00000a9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f000018f40000099c000012fc00003efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0011fff",
		x"f000014f4000009ac00001afc000016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009fff",
		x"f00000844000009b4000009cc00000d1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f000013f4000009dc000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f00003dfc00000f1c000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00b7fff",
		x"f00001dfc00000c9c000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0077fff",
		x"f00000844000009ec00000f14000009fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003bff",
		x"f000013f400000a0c00001ffc00009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f00000a8400000a1c00000e1c00000f1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00023ff",
		x"f00001ffc00000f1c00005ffc0000dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003ffff",
		x"f00000d0400000a2c0000121c00001a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00043ff",
		x"f0000140400000a3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a1",
		x"f00000ffc00000ebc0000117c0000197c00001efc00001efc000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000c00009ff",
		x"f00000ffc00000ebc0000157c00001d7c000013fc000013fc00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f000017fc0000137c00001bfc00001bfc000037fc000017fc0000dffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00001ffc00001b7c000017fc000017fc000037fc00001ffc0000bffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00000f7c00000c3c00000ebc00000ebc000013fc00001bfc00009ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000c0000dff",
		x"f00000cfc00000e3c00000fbc00000fbc00001bfc000017fc00003ffc0000bffb0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000efc00000fbc00001f7c000010fc000017fc000037fc0000fffc0001dffb0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000ffc00000fbc000018fc000014fc00001ffc00003ffc00001ffc00013ffb0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f00000ffc00000e7c00001cfc000012fc00001ffc00003ffc00009ffc0001bffb0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000ffc00000e7c00001afc000016fc000017fc000037fc00017ffc0000fffb0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00000abc00000ab400000a4400000a5c0000177c00003dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f00000db400000a6c00001fbc0000107c00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000fb400000a7c0000187c0000147c00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00011ff",
		x"f00000c7400000a8c00001c7c0000127c00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00009ff",
		x"f00000f7c00001a7c00001f7c00001f7c0000bffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002bff",
		x"f00000f7c0000167c000012fc000012fc0000fffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f00000e7400000a9c00001e7c0000117c000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00019ff",
		x"f00000efc0000197c00001afc00001afc00009ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003bff",
		x"f0000083c0000062400000aa400000abc000017fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000e7400000acc00000ddc00000fdc00003ffc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001dff",
		x"f00000efc00000c3c0000137c00001b7c0000fffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f00000efc00000e3c0000177c00001f7c00009ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f00000ff400000adc000010fc000018fc0000dffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000b7c000008d400000ae400000afc00001ffc00009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003bff",
		x"f000015fc00000f7c00001bfc00001bfc00027ffc00067ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00000afc0000083400000b0400000b1c00005ffc0000dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00001ffc000017fc000077fc00001ffc000dfffc001bfffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003ffff",
		x"f0000061400000b2c0000081400000b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f0000066400000b4400000b5400000b6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000e7400000b7c0000197c0000157b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00047ff",
		x"f00000e7400000b8c00001d7c00001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00000e7400000b9c0000137c000012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00067ff",
		x"f0000066400000bac00000b9c00000a5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00013ff",
		x"f00001cfc00000b5c000036fc000016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0019fff",
		x"f000012fc00000adc000036fc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00001afc00000bdc00003efc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0015fff",
		x"f000008c400000bb400000bcc00000e9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003bff",
		x"f000013f400000bdc00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0047fff",
		x"f00001bf400000bec00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0027fff",
		x"f000008c400000bfc00000c9400000c0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007bff",
		x"f000013f400000c1c00009ffc00019ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c009ffff",
		x"f00001bf400000c2c00005ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c005ffff",
		x"f00000b8400000c3c00000f1c00000f1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00063ff",
		x"f00000f0400000c4c0000161c00001e1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000c3ff",
		x"f00001c0400000c5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a1",
		x"f00000ef400000c6c000016fc000016fc0000dffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000efc0000157c00001efc00001efc0000bffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00000ef400000c7c000012fc000012fc0000fffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f00000ffc00001d7c00001afc00001afc00009ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f00000d7400000c8c000016fc000016fc0000dffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000ffc0000137c00001efc00001efc0000bffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000d7400000c9c00000fbc00000fbc000057fc000037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f00000f7400000cac00000e7c00000e7c000077fc0000bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00013ff",
		x"f00000cfc00000b5c00000e7c00000e7c000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f00001ffc00000f7c00001ffc00001ffc0001bffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f00001dfc00000f7c000017fc00001ffc00017ffc00057ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f000013fc00000efc00001ffc00003ffc00037ffc00077ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0017fff",
		x"f00001bfc00000efc000013fc000013fc0000fffc0004fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f000017fc00000efc00001bfc000017fc0002fffc0006fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f0000085400000cb400000cc400000cdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000ef400000ce400000cfc0000177b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f0000081400000d0400000d1c00000aeb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000f7400000d2c00001b7c000012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f000014fc00000bec00001afc00001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000f7400000d3c0000177c000016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00057ff",
		x"f00001cfc00000a1c000016fc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000afff",
		x"f000012fc00000b1c00001efc000012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f0000061400000d4c00000a3400000d5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f0000082400000d6400000d7c00000d9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00001bf400000d8c00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0067fff",
		x"f000017f400000d9c00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0017fff",
		x"f000017f400000dac000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0057fff",
		x"f0000082400000dbc00000e9c00000f5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00001ffc00000f5c0000dffc00015ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00dffff",
		x"f00003ffc00000f5c00003ffc0000dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00fffff",
		x"f00001bfc00000f5c0000bffc0001dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c01fffff",
		x"f00000a4400000dcc00000e9c00000e9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00013ff",
		x"f00000c8400000ddc0000111c0000191b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00023ff",
		x"f0000120400000deb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000161",
		x"f00001bfc000013fc00001dfc00003dfc00005ffc00015ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f000017fc000013fc000017fc000037fc0000dffc0001dffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00001ffc00001bfc000017fc000037fc00003ffc00013ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f00000ffc00000d3c000014fc00001cfc00007ffc0000fffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000ffc00000f3c000012fc00001afc00001ffc00009ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f000008d400000dfc00000a9c00000b9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000037f",
		x"f00000efc00000a5c00001f7c000010fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f000011fc00000b5c000018fc000014fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000efc00000adc00001cfc000012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00003ffc00001afc000077fc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f0000089400000e0c00000a9c00000b9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00000f7c00000a5c000012fc00001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00077ff",
		x"f00000f7c00000b5c00001afc000016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000efc00000adc000016fc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004fff",
		x"f0000065400000e1c00000b3400000e2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f000016f400000e3c00003efc000015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000dfff",
		x"f000008a400000e4400000e5c00000f9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00003df400000e6c000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00f7fff",
		x"f000017f400000e7c000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f000037f400000e8c000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c008ffff",
		x"f000017f400000e9c00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c004ffff",
		x"f00000aa400000eac00000d9c00000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00047ff",
		x"f00000b4400000ebc00000e9c00000e9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00053ff",
		x"f00000e8400000ecc0000151c00001d1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000a3ff",
		x"f00001a0400000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000161",
		x"f00000a3400000eec00000bd400000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f0000085400000f0c00000bd400000f1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00009ff",
		x"f0000083400000f2c00000ab400000f3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00001ef400000f4c000035fc000015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001dfff",
		x"f00001ef400000f5c000035fc00001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003dfff",
		x"f0000086400000f6400000f7c00000c5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f000037f400000f8c00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00cffff",
		x"f00001ffc00000e5c00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c002ffff",
		x"f00003ffc00000d5c00003ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00affff",
		x"f00001ffc00000f5c000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c006ffff",
		x"f00003ff400000f9c000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00effff",
		x"f00000ba400000fac00000f9c00000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00000ac400000fbc00000f9c00000f9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00033ff",
		x"f00000d8400000fcc0000131c00001b1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00063ff",
		x"f0000160400000fdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e1",
		x"f00000b3400000fe400000ff40000100b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f000019f40000101c00001efc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f000008d40000102c00000a340000103b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00005ff",
		x"f00001af40000104c00001efc000035fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006fff",
		x"f000008b400001054000010640000107b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f000013f40000108c00003dfc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f000013f40000109c00001dfc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0023fff",
		x"f00001bf4000010ac00003dfc000037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0013fff",
		x"f000008e4000010bc00000cdc00000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f000017fc00000ddc000017fc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f000037fc00000fdc000037fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c009ffff",
		x"f000017fc00000c3c00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c005ffff",
		x"f00000a64000010cc00000c5c00000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00067ff",
		x"f00000bc4000010dc00000f9c00000f9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00073ff",
		x"f00000f84000010ec0000171c00001f1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000e3ff",
		x"f00001e04000010fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e1",
		x"f00000ab40000110c00000c3c00000e3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f000015f40000111c000013fc000013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f00001dfc00000d3c00001bfc00001bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006fff",
		x"f000013fc00000f3c000017fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f0000083400001124000011340000114b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000dff",
		x"f000016f40000115c000013fc000015fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000efff",
		x"f00001ef40000116c000013fc000035fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f0000087c00000204000011740000118b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00001bf40000119c000015fc000035fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0033fff",
		x"f000017f4000011ac000015fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000bfff",
		x"f000017fc00000dbc000035fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c002bfff",
		x"f00001ffc00000fbc00001dfc000057fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001bfff",
		x"f00001ffc00000c7c00003dfc000037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003bfff",
		x"f00000814000011bc00000e3c00000d3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00077ff",
		x"f00000b64000011cc00000e5c00000edb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f00000a24000011dc00000e5c00000e5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f00000c44000011ec0000109c0000189b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00013ff",
		x"f00001104000011fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000121",
		x"f00000bbc0000060c00000cb40000120b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000dff",
		x"f00001bfc00000ebc00001ffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00000ab4000012140000122c00000d3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00003ff",
		x"f000011f40000123c00001bfc00001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009fff",
		x"f000019fc00000f3c00003dfc00001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f000015fc00000cbc00003dfc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00001dfc00000ebc000037fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000dfff",
		x"f000013f40000124c00001dfc00003dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f000013fc00000e7c000017fc000077fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0027fff",
		x"f00001bf40000125c000037fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0017fff",
		x"f00001bfc00000d7c000037fc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0037fff",
		x"f000008940000126c00000f3c00000cbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000ae4000012740000128c00000fdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00057ff",
		x"f00000b240000129c00000e5c0000113b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004bff",
		x"f00000e44000012ac0000149c00001c9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00093ff",
		x"f00001904000012bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000121",
		x"f000017f4000012cc00003ffc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00000bbc00000404000012dc00000dbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f000013f4000012ec000037fc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00001bf4000012fc00001bfc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000bfff",
		x"f000017f40000130c00001ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f000017f40000131c00003ffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c002ffff",
		x"f000008540000132c00000ebc00000dbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004fff",
		x"f00000be4000013340000134c00000fdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f000017f40000135c00007ffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003ffff",
		x"f00000aa40000136c00000e5c0000193b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002bff",
		x"f00000d440000137c0000129c00001a9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00053ff",
		x"f000015040000138b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a1",
		x"f00001ffc00000f7c000037fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00001ffc00000fbc00001ffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0017fff",
		x"f00001ffc00000c7c000017fc000037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f000017fc00000e7c000017fc000037fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f00001ffc00000f7c00001ffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f00001ffc00000cfc00003ffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003ffff",
		x"f000008d40000139c00000fb4000013ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000a14000013bc00000fdc00000fdb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00077ff",
		x"f000017fc00000e3c0000fffc00013ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00bffff",
		x"f00001ffc00000e3c00001ffc0000bffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c007ffff",
		x"f00000ba4000013cc00000f5c0000153b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006bff",
		x"f00000f44000013dc0000169c00001e9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000d3ff",
		x"f00001d04000013eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a1",
		x"f00000834000013fc00000c740000140b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006fff",
		x"f000037f40000141c0000dffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00dffff",
		x"f00000b140000142c00000e3c00000e3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000a640000143c00000f5c00001d3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f00000cc40000144c0000119c0000199b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00033ff",
		x"f000013040000145b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000161",
		x"f000008b40000146c00000e740000147b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00001ffc00000efc0000bffc00007ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c003ffff",
		x"f00003ff40000148c0000fffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00bffff",
		x"f00000a940000149c00000f3c00000f3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004fff",
		x"f00000b64000014ac00000f5c0000133b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005bff",
		x"f00000ec4000014bc0000159c00001d9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000b3ff",
		x"f00001b04000014cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000161",
		x"f00000874000014dc00000d7c00000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00001ffc00000efc00009ffc00005ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c007ffff",
		x"f00003ffc00000efc0000dffc00003ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00fffff",
		x"f00000b94000014ec00000f3c00000f3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000cfff",
		x"f00000ae4000014fc00000f5c00001b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003bff",
		x"f00000dc40000150c0000139c00001b9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00073ff",
		x"f000017040000151b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e1",
		x"f00000afc0000020c00000f7c00000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00000a540000152c00000ebc00000ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000be40000153c00000edc0000173b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007bff",
		x"f00000fc40000154c0000179c00001f9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000f3ff",
		x"f00001f040000155b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e1",
		x"f00000b540000156c00000ebc00000ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000afff",
		x"f00000a140000157c00000edc00001f3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f00000c240000158c0000105c0000185b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000bff",
		x"f000010840000159b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000131",
		x"f00000ad4000015ac00000fbc00000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006fff",
		x"f00000b14000015bc00000edc000010bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00047ff",
		x"f00000e24000015cc0000145c00001c5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0008bff",
		x"f00001884000015db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000131",
		x"f00000bd4000015ec00000fbc00000fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000efff",
		x"f00000c94000015fc00000edc000018bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00000d240000160c0000125c00001a5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004bff",
		x"f000014840000161b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b1",
		x"f00000a340000162c00000e7c00000e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00000e940000163c00000fdc000014bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000a7ff",
		x"f00000f240000164c0000165c00001e5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000cbff",
		x"f00001c840000165b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b1",
		x"f00000b340000166c00000e7c00000e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009fff",
		x"f00000d940000167c00000fdc00001cbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00067ff",
		x"f00000ca40000168c0000115c0000195b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002bff",
		x"f000012840000169b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000171",
		x"f00000ab4000016ac00000f7c00000f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00000f94000016bc00000fdc000012bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000e7ff",
		x"f00000ea4000016cc0000155c000016bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000abff",
		x"f00001a84000016db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000171",
		x"f00000bb4000016ec00000f7c00000f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000dfff",
		x"f00000c54000016fc00000fdc00001abb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f00000da40000170c00001d5c000016bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006bff",
		x"f000016840000171b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f1",
		x"f00000a740000172c00000efc00000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00000e540000173c00000e3c000016bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00097ff",
		x"f00000fa40000174c0000135c00001ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ebff",
		x"f00001e840000175b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f1",
		x"f00000b740000176c00000efc00000efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000bfff",
		x"f00000d540000177c00000e3c00001ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00057ff",
		x"f00000c640000178c00001b5c00001ebb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001bff",
		x"f000011840000179b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000131",
		x"f00000af4000017ac00000ffc00000ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f00000f54000017bc00000e3c000011bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000d7ff",
		x"f00000e64000017cc0000175c000013bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009bff",
		x"f00001984000017db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000131",
		x"f00000dfc0000020c00000ffc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f00000cd4000017ec00000e3c000019bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f00000d64000017fc00001f5c000013bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005bff",
		x"f000015840000180b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b1",
		x"f00000ed40000181c000015bc00001dbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000b7ff",
		x"f00000f640000182c000010dc00001bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000dbff",
		x"f00001d840000183b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b1",
		x"f00000dd40000184c000013bc00001bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00077ff",
		x"f00000ce40000185c000018dc00001bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003bff",
		x"f000013840000186b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000171",
		x"f00000fd40000187c000017bc00001fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000f7ff",
		x"f00000ee40000188c000014dc000017bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000bbff",
		x"f00001b840000189b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000171",
		x"f00000c34000018ac0000107c0000187b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00000de4000018bc00001cdc000017bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007bff",
		x"f00001784000018cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f1",
		x"f00000e34000018dc0000147c00001c7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0008fff",
		x"f00000fe4000018ec000012dc00001fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000fbff",
		x"f00001f84000018fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f1",
		x"f00000d340000190c0000127c00001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004fff",
		x"f00000c140000191c00001adc00001fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00007ff",
		x"f000010440000192b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000129",
		x"f00000f340000193c0000167c00001e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000cfff",
		x"f00000e140000194c000016dc000013bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00087ff",
		x"f000018440000195b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000129",
		x"f00000cb40000196c0000117c0000197b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00000d140000197c00001edc000013bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00047ff",
		x"f000014440000198b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a9",
		x"f00000eb40000199c0000157c00001d7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000afff",
		x"f00000f14000019ac000011dc00001bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000c7ff",
		x"f00001c44000019bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a9",
		x"f00000db4000019cc0000137c00001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006fff",
		x"f00000c94000019dc000019dc00001bbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00027ff",
		x"f00001244000019eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000169",
		x"f00000fb4000019fc0000177c00001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000efff",
		x"f00000e9400001a0c000015dc000017bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000a7ff",
		x"f00001a4400001a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000169",
		x"f00000c7400001a2c000010fc000018fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00000d9400001a3c00001ddc000017bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00067ff",
		x"f0000164400001a4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e9",
		x"f00000e7400001a5c000014fc00001cfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009fff",
		x"f00000f9400001a6c000013dc00001fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000e7ff",
		x"f00001e4400001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e9",
		x"f00000d7400001a8c000012fc00001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f00000c5400001a9c00001bdc00001fbb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00017ff",
		x"f0000114400001aab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000129",
		x"f00000f7400001abc000016fc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000dfff",
		x"f00000e5400001acc000017dc0000127b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00097ff",
		x"f0000194400001adb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000129",
		x"f00000cf400001aec000011fc000019fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00000d5400001afc00001fdc0000127b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00057ff",
		x"f0000154400001b0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a9",
		x"f00000ef400001b1c000015fc00001dfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000bfff",
		x"f00000f5400001b2c0000103c00001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000d7ff",
		x"f00001d4400001b3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a9",
		x"f00000df400001b4c000013fc00001bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f00000f5400001b5c0000183c00001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001d7ff",
		x"f0000134400001b6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000169",
		x"f00000ffc0000020c000017fc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f00000ed400001b7c0000143c0000167b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00037ff",
		x"f00001b4400001b8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000169",
		x"f00000ed400001b9c00001c3c0000167b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00137ff",
		x"f0000174400001bab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e9",
		x"f00000ed400001bbc0000123c00001e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000b7ff",
		x"f00001f4400001bcb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e9",
		x"f00000ed400001bdc00001a3c00001e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001b7ff",
		x"f000010c400001beb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000139",
		x"f00000fd400001bfc0000163c0000127b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00077ff",
		x"f000018c400001c0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000139",
		x"f00000fd400001c1c00001e3c0000127b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00177ff",
		x"f000014c400001c2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b9",
		x"f00000fd400001c3c0000113c00001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000f7ff",
		x"f00001cc400001c4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b9",
		x"f00000fd400001c5c0000193c00001a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001f7ff",
		x"f000012c400001c6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000179",
		x"f00000e3400001c7c0000153c0000167b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000fff",
		x"f00001ac400001c8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000179",
		x"f00000e3400001c9c00001d3c0000167b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0010fff",
		x"f000016c400001cab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f9",
		x"f00000e3400001cbc0000133c00001e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0008fff",
		x"f00001ec400001ccb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f9",
		x"f00000e3400001cdc00001b3c00001e7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0018fff",
		x"f000011c400001ceb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000139",
		x"f00000f3400001cfc0000173c0000137b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0004fff",
		x"f000019c400001d0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000139",
		x"f00000f3400001d1c00001f3c0000137b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0014fff",
		x"f000015c400001d2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b9",
		x"f00000f3400001d3c000010bc00001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000cfff",
		x"f00001dc400001d4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b9",
		x"f00000f3400001d5c000018bc00001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001cfff",
		x"f000013c400001d6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000179",
		x"f00000eb400001d7c000014bc0000177b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0002fff",
		x"f00001bc400001d8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000179",
		x"f00000eb400001d9c00001cbc0000177b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0012fff",
		x"f000017c400001dab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f9",
		x"f00000eb400001dbc000012bc00001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000afff",
		x"f00001fc400001dcb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f9",
		x"f00000eb400001ddc00001abc00001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001afff",
		x"f0000102400001deb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000125",
		x"f00000fb400001dfc0000137c0000137b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0006fff",
		x"f0000182400001e0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000125",
		x"f00000fb400001e1c00001b7c00001b7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0016fff",
		x"f0000142400001e2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a5",
		x"f00000fb400001e3c0000177c0000177b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000efff",
		x"f00001c2400001e4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a5",
		x"f00000fb400001e5c00001f7c00001f7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001efff",
		x"f0000122400001e6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000165",
		x"f00000e7400001e7c000012fc000012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0001fff",
		x"f00001a2400001e8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000165",
		x"f00000e7400001e9c00001afc00001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0011fff",
		x"f0000162400001eab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e5",
		x"f00000e7400001ebc000016fc000016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0009fff",
		x"f00001e2400001ecb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e5",
		x"f00000e7400001edc00001efc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0019fff",
		x"f0000112400001eeb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000125",
		x"f00000f7400001efc000012fc000012fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0005fff",
		x"f0000192400001f0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000125",
		x"f00000f7400001f1c00001afc00001afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0015fff",
		x"f0000152400001f2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a5",
		x"f00000f7400001f3c000016fc000016fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000dfff",
		x"f00001d2400001f4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a5",
		x"f00000f7400001f5c00001efc00001efb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001dfff",
		x"f0000132400001f6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000165",
		x"f00000ef400001f7c000013fc000013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0003fff",
		x"f00001b2400001f8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000165",
		x"f00000ef400001f9c00001bfc00001bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0013fff",
		x"f0000172400001fab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e5",
		x"f00000ef400001fbc000017fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000bfff",
		x"f00001f2400001fcb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e5",
		x"f00000ef400001fdc00001ffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001bfff",
		x"f000010a400001feb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000135",
		x"f00000ff400001ffc000013fc000013fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0007fff",
		x"f000018a40000200b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000135",
		x"f00000ff40000201c00001bfc00001bfb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0017fff",
		x"f000014a40000202b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b5",
		x"f00000ff40000203c000017fc000017fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000ffff",
		x"f00001ca40000204b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b5",
		x"f00000ffc0000020c00001ffc00001ffb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c001ffff",
		x"f000012a40000205b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000175",
		x"f00001aa40000206b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000175",
		x"f000016a40000207b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f5",
		x"f00001ea40000208b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f5",
		x"f000011a40000209b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000135",
		x"f000019a4000020ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000135",
		x"f000015a4000020bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b5",
		x"f00001da4000020cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b5",
		x"f000013a4000020db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000175",
		x"f00001ba4000020eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000175",
		x"f000017a4000020fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f5",
		x"f00001fa40000210b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f5",
		x"f000010640000211b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012d",
		x"f000018640000212b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012d",
		x"f000014640000213b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ad",
		x"f00001c640000214b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ad",
		x"f000012640000215b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016d",
		x"f00001a640000216b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016d",
		x"f000016640000217b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ed",
		x"f00001e640000218b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ed",
		x"f000011640000219b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012d",
		x"f00001964000021ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012d",
		x"f00001564000021bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ad",
		x"f00001d64000021cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ad",
		x"f00001364000021db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016d",
		x"f00001b64000021eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016d",
		x"f00001764000021fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ed",
		x"f00001f640000220b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ed",
		x"f000010e40000221b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013d",
		x"f000018e40000222b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013d",
		x"f000014e40000223b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bd",
		x"f00001ce40000224b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bd",
		x"f000012e40000225b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017d",
		x"f00001ae40000226b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017d",
		x"f000016e40000227b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fd",
		x"f00001ee40000228b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fd",
		x"f000011e40000229b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013d",
		x"f000019e4000022ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013d",
		x"f000015e4000022bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bd",
		x"f00001de4000022cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bd",
		x"f000013e4000022db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017d",
		x"f00001be4000022eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017d",
		x"f000017e4000022fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fd",
		x"f00001fe40000230b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fd",
		x"f000010140000231b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000123",
		x"f000018140000232b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000123",
		x"f000014140000233b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a3",
		x"f00001c140000234b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a3",
		x"f000012140000235b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000163",
		x"f00001a140000236b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000163",
		x"f000016140000237b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e3",
		x"f00001e140000238b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e3",
		x"f000011140000239b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000123",
		x"f00001914000023ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000123",
		x"f00001514000023bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a3",
		x"f00001d14000023cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a3",
		x"f00001314000023db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000163",
		x"f00001b14000023eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000163",
		x"f00001714000023fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e3",
		x"f00001f140000240b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e3",
		x"f000010940000241b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000133",
		x"f000018940000242b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000133",
		x"f000014940000243b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b3",
		x"f00001c940000244b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b3",
		x"f000012940000245b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000173",
		x"f00001a940000246b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000173",
		x"f000016940000247b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f3",
		x"f00001e940000248b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f3",
		x"f000011940000249b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000133",
		x"f00001994000024ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000133",
		x"f00001594000024bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b3",
		x"f00001d94000024cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b3",
		x"f00001394000024db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000173",
		x"f00001b94000024eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000173",
		x"f00001794000024fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f3",
		x"f00001f940000250b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f3",
		x"f000010540000251b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012b",
		x"f000018540000252b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012b",
		x"f000014540000253b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ab",
		x"f00001c540000254b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ab",
		x"f000012540000255b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016b",
		x"f00001a540000256b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016b",
		x"f000016540000257b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001eb",
		x"f00001e540000258b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001eb",
		x"f000011540000259b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012b",
		x"f00001954000025ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012b",
		x"f00001554000025bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ab",
		x"f00001d54000025cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ab",
		x"f00001354000025db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016b",
		x"f00001b54000025eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016b",
		x"f00001754000025fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001eb",
		x"f00001f540000260b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001eb",
		x"f000010d40000261b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013b",
		x"f000018d40000262b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013b",
		x"f000014d40000263b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bb",
		x"f00001cd40000264b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bb",
		x"f000012d40000265b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017b",
		x"f00001ad40000266b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017b",
		x"f000016d40000267b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fb",
		x"f00001ed40000268b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fb",
		x"f000011d40000269b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013b",
		x"f000019d4000026ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013b",
		x"f000015d4000026bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bb",
		x"f00001dd4000026cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bb",
		x"f000013d4000026db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017b",
		x"f00001bd4000026eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017b",
		x"f000017d4000026fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fb",
		x"f00001fd40000270b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001fb",
		x"f000010340000271b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000127",
		x"f000018340000272b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000127",
		x"f000014340000273b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a7",
		x"f00001c340000274b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a7",
		x"f000012340000275b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000167",
		x"f00001a340000276b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000167",
		x"f000016340000277b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e7",
		x"f00001e340000278b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e7",
		x"f000011340000279b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000127",
		x"f00001934000027ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000127",
		x"f00001534000027bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a7",
		x"f00001d34000027cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001a7",
		x"f00001334000027db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000167",
		x"f00001b34000027eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000167",
		x"f00001734000027fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e7",
		x"f00001f340000280b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001e7",
		x"f000010b40000281b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000137",
		x"f000018b40000282b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000137",
		x"f000014b40000283b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b7",
		x"f00001cb40000284b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b7",
		x"f000012b40000285b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000177",
		x"f00001ab40000286b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000177",
		x"f000016b40000287b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f7",
		x"f00001eb40000288b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f7",
		x"f000011b40000289b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000137",
		x"f000019b4000028ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000137",
		x"f000015b4000028bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b7",
		x"f00001db4000028cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001b7",
		x"f000013b4000028db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000177",
		x"f00001bb4000028eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c0000177",
		x"f000017b4000028fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f7",
		x"f00001fb40000290b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001f7",
		x"f000010740000291b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012f",
		x"f000018740000292b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012f",
		x"f000014740000293b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001af",
		x"f00001c740000294b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001af",
		x"f000012740000295b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00001a740000296b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f000016740000297b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ef",
		x"f00001e740000298b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ef",
		x"f000011740000299b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012f",
		x"f00001974000029ab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000012f",
		x"f00001574000029bb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001af",
		x"f00001d74000029cb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001af",
		x"f00001374000029db0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00001b74000029eb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000016f",
		x"f00001774000029fb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ef",
		x"f00001f7400002a0b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ef",
		x"f000010f400002a1b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013f",
		x"f000018f400002a2b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013f",
		x"f000014f400002a3b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bf",
		x"f00001cf400002a4b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bf",
		x"f000012f400002a5b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f00001af400002a6b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f000016f400002a7b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00001ef400002a8b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f000011f400002a9b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013f",
		x"f000019f400002aab0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000013f",
		x"f000015f400002abb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bf",
		x"f00001df400002acb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001bf",
		x"f000013f400002adb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f00001bf400002aeb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c000017f",
		x"f000017f400002afb0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff",
		x"f00001ffc0000020b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000b0000000c00001ff"
    );
end ccsds_constants;

package body ccsds_constants is
	
end ccsds_constants;
